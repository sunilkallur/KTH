
module SRAM ( rst_n, rws, addrs, inp, outp );
  input [2:0] addrs;
  input [15:0] inp;
  output [15:0] outp;
  input rst_n, rws;
  wire   \mem2[0][15] , \mem2[0][14] , \mem2[0][13] , \mem2[0][12] ,
         \mem2[0][11] , \mem2[0][10] , \mem2[0][9] , \mem2[0][8] ,
         \mem2[0][7] , \mem2[0][6] , \mem2[0][5] , \mem2[0][4] , \mem2[0][3] ,
         \mem2[0][2] , \mem2[0][1] , \mem2[0][0] , \mem2[1][15] ,
         \mem2[1][14] , \mem2[1][13] , \mem2[1][12] , \mem2[1][11] ,
         \mem2[1][10] , \mem2[1][9] , \mem2[1][8] , \mem2[1][7] , \mem2[1][6] ,
         \mem2[1][5] , \mem2[1][4] , \mem2[1][3] , \mem2[1][2] , \mem2[1][1] ,
         \mem2[1][0] , \mem2[2][15] , \mem2[2][14] , \mem2[2][13] ,
         \mem2[2][12] , \mem2[2][11] , \mem2[2][10] , \mem2[2][9] ,
         \mem2[2][8] , \mem2[2][7] , \mem2[2][6] , \mem2[2][5] , \mem2[2][4] ,
         \mem2[2][3] , \mem2[2][2] , \mem2[2][1] , \mem2[2][0] , \mem2[3][15] ,
         \mem2[3][14] , \mem2[3][13] , \mem2[3][12] , \mem2[3][11] ,
         \mem2[3][10] , \mem2[3][9] , \mem2[3][8] , \mem2[3][7] , \mem2[3][6] ,
         \mem2[3][5] , \mem2[3][4] , \mem2[3][3] , \mem2[3][2] , \mem2[3][1] ,
         \mem2[3][0] , \mem2[4][15] , \mem2[4][14] , \mem2[4][13] ,
         \mem2[4][12] , \mem2[4][11] , \mem2[4][10] , \mem2[4][9] ,
         \mem2[4][8] , \mem2[4][7] , \mem2[4][6] , \mem2[4][5] , \mem2[4][4] ,
         \mem2[4][3] , \mem2[4][2] , \mem2[4][1] , \mem2[4][0] , N47, N48, N49,
         N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63,
         N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77,
         N78, N79, N80, N81, N82, N83, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n1, n2, n3, n4, n5, n49, n50, n51, n52,
         n53, n54, n55, n56;

  LHD1 \mem2_reg[0][15]  ( .E(N66), .D(N62), .Q(\mem2[0][15] ) );
  LHD1 \mem2_reg[0][14]  ( .E(N66), .D(N61), .Q(\mem2[0][14] ) );
  LHD1 \mem2_reg[0][13]  ( .E(N66), .D(N60), .Q(\mem2[0][13] ) );
  LHD1 \mem2_reg[0][12]  ( .E(N66), .D(N59), .Q(\mem2[0][12] ) );
  LHD1 \mem2_reg[0][11]  ( .E(N66), .D(N58), .Q(\mem2[0][11] ) );
  LHD1 \mem2_reg[0][10]  ( .E(N66), .D(N57), .Q(\mem2[0][10] ) );
  LHD1 \mem2_reg[0][9]  ( .E(N66), .D(N56), .Q(\mem2[0][9] ) );
  LHD1 \mem2_reg[0][8]  ( .E(N66), .D(N55), .Q(\mem2[0][8] ) );
  LHD1 \mem2_reg[0][7]  ( .E(N66), .D(N54), .Q(\mem2[0][7] ) );
  LHD1 \mem2_reg[0][6]  ( .E(N66), .D(N53), .Q(\mem2[0][6] ) );
  LHD1 \mem2_reg[0][5]  ( .E(N66), .D(N52), .Q(\mem2[0][5] ) );
  LHD1 \mem2_reg[0][4]  ( .E(N66), .D(N51), .Q(\mem2[0][4] ) );
  LHD1 \mem2_reg[0][3]  ( .E(N66), .D(N50), .Q(\mem2[0][3] ) );
  LHD1 \mem2_reg[0][2]  ( .E(N66), .D(N49), .Q(\mem2[0][2] ) );
  LHD1 \mem2_reg[0][1]  ( .E(N66), .D(N48), .Q(\mem2[0][1] ) );
  LHD1 \mem2_reg[0][0]  ( .E(N66), .D(N47), .Q(\mem2[0][0] ) );
  LHD1 \mem2_reg[1][15]  ( .E(N65), .D(N62), .Q(\mem2[1][15] ) );
  LHD1 \mem2_reg[1][14]  ( .E(N65), .D(N61), .Q(\mem2[1][14] ) );
  LHD1 \mem2_reg[1][13]  ( .E(N65), .D(N60), .Q(\mem2[1][13] ) );
  LHD1 \mem2_reg[1][12]  ( .E(N65), .D(N59), .Q(\mem2[1][12] ) );
  LHD1 \mem2_reg[1][11]  ( .E(N65), .D(N58), .Q(\mem2[1][11] ) );
  LHD1 \mem2_reg[1][10]  ( .E(N65), .D(N57), .Q(\mem2[1][10] ) );
  LHD1 \mem2_reg[1][9]  ( .E(N65), .D(N56), .Q(\mem2[1][9] ) );
  LHD1 \mem2_reg[1][8]  ( .E(N65), .D(N55), .Q(\mem2[1][8] ) );
  LHD1 \mem2_reg[1][7]  ( .E(N65), .D(N54), .Q(\mem2[1][7] ) );
  LHD1 \mem2_reg[1][6]  ( .E(N65), .D(N53), .Q(\mem2[1][6] ) );
  LHD1 \mem2_reg[1][5]  ( .E(N65), .D(N52), .Q(\mem2[1][5] ) );
  LHD1 \mem2_reg[1][4]  ( .E(N65), .D(N51), .Q(\mem2[1][4] ) );
  LHD1 \mem2_reg[1][3]  ( .E(N65), .D(N50), .Q(\mem2[1][3] ) );
  LHD1 \mem2_reg[1][2]  ( .E(N65), .D(N49), .Q(\mem2[1][2] ) );
  LHD1 \mem2_reg[1][1]  ( .E(N65), .D(N48), .Q(\mem2[1][1] ) );
  LHD1 \mem2_reg[1][0]  ( .E(N65), .D(N47), .Q(\mem2[1][0] ) );
  LHD1 \mem2_reg[2][15]  ( .E(N64), .D(N62), .Q(\mem2[2][15] ) );
  LHD1 \mem2_reg[2][14]  ( .E(N64), .D(N61), .Q(\mem2[2][14] ) );
  LHD1 \mem2_reg[2][13]  ( .E(N64), .D(N60), .Q(\mem2[2][13] ) );
  LHD1 \mem2_reg[2][12]  ( .E(N64), .D(N59), .Q(\mem2[2][12] ) );
  LHD1 \mem2_reg[2][11]  ( .E(N64), .D(N58), .Q(\mem2[2][11] ) );
  LHD1 \mem2_reg[2][10]  ( .E(N64), .D(N57), .Q(\mem2[2][10] ) );
  LHD1 \mem2_reg[2][9]  ( .E(N64), .D(N56), .Q(\mem2[2][9] ) );
  LHD1 \mem2_reg[2][8]  ( .E(N64), .D(N55), .Q(\mem2[2][8] ) );
  LHD1 \mem2_reg[2][7]  ( .E(N64), .D(N54), .Q(\mem2[2][7] ) );
  LHD1 \mem2_reg[2][6]  ( .E(N64), .D(N53), .Q(\mem2[2][6] ) );
  LHD1 \mem2_reg[2][5]  ( .E(N64), .D(N52), .Q(\mem2[2][5] ) );
  LHD1 \mem2_reg[2][4]  ( .E(N64), .D(N51), .Q(\mem2[2][4] ) );
  LHD1 \mem2_reg[2][3]  ( .E(N64), .D(N50), .Q(\mem2[2][3] ) );
  LHD1 \mem2_reg[2][2]  ( .E(N64), .D(N49), .Q(\mem2[2][2] ) );
  LHD1 \mem2_reg[2][1]  ( .E(N64), .D(N48), .Q(\mem2[2][1] ) );
  LHD1 \mem2_reg[2][0]  ( .E(N64), .D(N47), .Q(\mem2[2][0] ) );
  LHD1 \mem2_reg[3][15]  ( .E(N63), .D(N62), .Q(\mem2[3][15] ) );
  LHD1 \mem2_reg[3][14]  ( .E(N63), .D(N61), .Q(\mem2[3][14] ) );
  LHD1 \mem2_reg[3][13]  ( .E(N63), .D(N60), .Q(\mem2[3][13] ) );
  LHD1 \mem2_reg[3][12]  ( .E(N63), .D(N59), .Q(\mem2[3][12] ) );
  LHD1 \mem2_reg[3][11]  ( .E(N63), .D(N58), .Q(\mem2[3][11] ) );
  LHD1 \mem2_reg[3][10]  ( .E(N63), .D(N57), .Q(\mem2[3][10] ) );
  LHD1 \mem2_reg[3][9]  ( .E(N63), .D(N56), .Q(\mem2[3][9] ) );
  LHD1 \mem2_reg[3][8]  ( .E(N63), .D(N55), .Q(\mem2[3][8] ) );
  LHD1 \mem2_reg[3][7]  ( .E(N63), .D(N54), .Q(\mem2[3][7] ) );
  LHD1 \mem2_reg[3][6]  ( .E(N63), .D(N53), .Q(\mem2[3][6] ) );
  LHD1 \mem2_reg[3][5]  ( .E(N63), .D(N52), .Q(\mem2[3][5] ) );
  LHD1 \mem2_reg[3][4]  ( .E(N63), .D(N51), .Q(\mem2[3][4] ) );
  LHD1 \mem2_reg[3][3]  ( .E(N63), .D(N50), .Q(\mem2[3][3] ) );
  LHD1 \mem2_reg[3][2]  ( .E(N63), .D(N49), .Q(\mem2[3][2] ) );
  LHD1 \mem2_reg[3][1]  ( .E(N63), .D(N48), .Q(\mem2[3][1] ) );
  LHD1 \mem2_reg[3][0]  ( .E(N63), .D(N47), .Q(\mem2[3][0] ) );
  LNCND1 \mem2_reg[4][15]  ( .D(inp[15]), .EN(n48), .CDN(rst_n), .Q(
        \mem2[4][15] ) );
  LNCND1 \mem2_reg[4][14]  ( .D(inp[14]), .EN(n48), .CDN(rst_n), .Q(
        \mem2[4][14] ) );
  LNCND1 \mem2_reg[4][13]  ( .D(inp[13]), .EN(n48), .CDN(rst_n), .Q(
        \mem2[4][13] ) );
  LNCND1 \mem2_reg[4][12]  ( .D(inp[12]), .EN(n48), .CDN(rst_n), .Q(
        \mem2[4][12] ) );
  LNCND1 \mem2_reg[4][11]  ( .D(inp[11]), .EN(n48), .CDN(rst_n), .Q(
        \mem2[4][11] ) );
  LNCND1 \mem2_reg[4][10]  ( .D(inp[10]), .EN(n48), .CDN(rst_n), .Q(
        \mem2[4][10] ) );
  LNCND1 \mem2_reg[4][9]  ( .D(inp[9]), .EN(n48), .CDN(rst_n), .Q(\mem2[4][9] ) );
  LNCND1 \mem2_reg[4][8]  ( .D(inp[8]), .EN(n48), .CDN(rst_n), .Q(\mem2[4][8] ) );
  LNCND1 \mem2_reg[4][7]  ( .D(inp[7]), .EN(n48), .CDN(rst_n), .Q(\mem2[4][7] ) );
  LNCND1 \mem2_reg[4][6]  ( .D(inp[6]), .EN(n48), .CDN(rst_n), .Q(\mem2[4][6] ) );
  LNCND1 \mem2_reg[4][5]  ( .D(inp[5]), .EN(n48), .CDN(rst_n), .Q(\mem2[4][5] ) );
  LNCND1 \mem2_reg[4][4]  ( .D(inp[4]), .EN(n48), .CDN(rst_n), .Q(\mem2[4][4] ) );
  LNCND1 \mem2_reg[4][3]  ( .D(inp[3]), .EN(n48), .CDN(rst_n), .Q(\mem2[4][3] ) );
  LNCND1 \mem2_reg[4][2]  ( .D(inp[2]), .EN(n48), .CDN(rst_n), .Q(\mem2[4][2] ) );
  LNCND1 \mem2_reg[4][1]  ( .D(inp[1]), .EN(n48), .CDN(rst_n), .Q(\mem2[4][1] ) );
  LNCND1 \mem2_reg[4][0]  ( .D(inp[0]), .EN(n48), .CDN(rst_n), .Q(\mem2[4][0] ) );
  LHD1 \outp_reg[15]  ( .E(N67), .D(N83), .Q(outp[15]) );
  LHD1 \outp_reg[14]  ( .E(N67), .D(N82), .Q(outp[14]) );
  LHD1 \outp_reg[13]  ( .E(N67), .D(N81), .Q(outp[13]) );
  LHD1 \outp_reg[12]  ( .E(N67), .D(N80), .Q(outp[12]) );
  LHD1 \outp_reg[11]  ( .E(N67), .D(N79), .Q(outp[11]) );
  LHD1 \outp_reg[10]  ( .E(N67), .D(N78), .Q(outp[10]) );
  LHD1 \outp_reg[9]  ( .E(N67), .D(N77), .Q(outp[9]) );
  LHD1 \outp_reg[8]  ( .E(N67), .D(N76), .Q(outp[8]) );
  LHD1 \outp_reg[7]  ( .E(N67), .D(N75), .Q(outp[7]) );
  LHD1 \outp_reg[6]  ( .E(N67), .D(N74), .Q(outp[6]) );
  LHD1 \outp_reg[5]  ( .E(N67), .D(N73), .Q(outp[5]) );
  LHD1 \outp_reg[4]  ( .E(N67), .D(N72), .Q(outp[4]) );
  LHD1 \outp_reg[3]  ( .E(N67), .D(N71), .Q(outp[3]) );
  LHD1 \outp_reg[2]  ( .E(N67), .D(N70), .Q(outp[2]) );
  LHD1 \outp_reg[1]  ( .E(N67), .D(N69), .Q(outp[1]) );
  LHD1 \outp_reg[0]  ( .E(N67), .D(N68), .Q(outp[0]) );
  BUFFD0 U3 ( .I(n52), .Z(n49) );
  BUFFD0 U4 ( .I(n52), .Z(n50) );
  BUFFD0 U5 ( .I(n9), .Z(n4) );
  NR2D1 U6 ( .A1(n51), .A2(n44), .ZN(n9) );
  BUFFD0 U7 ( .I(n52), .Z(n51) );
  OAI21D1 U8 ( .A1(n43), .A2(n47), .B(rst_n), .ZN(N63) );
  OAI21D1 U9 ( .A1(n45), .A2(n47), .B(rst_n), .ZN(N64) );
  OAI21D1 U10 ( .A1(n46), .A2(n47), .B(rst_n), .ZN(N65) );
  ND2D1 U11 ( .A1(rst_n), .A2(n53), .ZN(N67) );
  ND3D1 U12 ( .A1(n55), .A2(n54), .A3(n56), .ZN(n44) );
  ND2D1 U13 ( .A1(n54), .A2(n53), .ZN(n47) );
  BUFFD0 U14 ( .I(n8), .Z(n3) );
  NR2D1 U15 ( .A1(n45), .A2(n49), .ZN(n8) );
  BUFFD0 U16 ( .I(n11), .Z(n1) );
  NR2D1 U17 ( .A1(n46), .A2(n49), .ZN(n11) );
  BUFFD0 U18 ( .I(n12), .Z(n2) );
  NR2D1 U19 ( .A1(n54), .A2(n50), .ZN(n12) );
  BUFFD0 U20 ( .I(n10), .Z(n5) );
  NR2D1 U21 ( .A1(n43), .A2(n50), .ZN(n10) );
  INVD1 U22 ( .I(rst_n), .ZN(n52) );
  OAI21D1 U23 ( .A1(rws), .A2(n44), .B(rst_n), .ZN(N66) );
  ND4D1 U24 ( .A1(addrs[2]), .A2(n56), .A3(n55), .A4(n53), .ZN(n48) );
  INVD1 U25 ( .I(addrs[2]), .ZN(n54) );
  ND2D1 U26 ( .A1(addrs[0]), .A2(n55), .ZN(n46) );
  ND2D1 U27 ( .A1(addrs[1]), .A2(n56), .ZN(n45) );
  ND2D1 U28 ( .A1(addrs[1]), .A2(addrs[0]), .ZN(n43) );
  INVD1 U29 ( .I(addrs[0]), .ZN(n56) );
  INVD1 U30 ( .I(rws), .ZN(n53) );
  INVD1 U31 ( .I(addrs[1]), .ZN(n55) );
  AN2D0 U32 ( .A1(inp[0]), .A2(rst_n), .Z(N47) );
  AN2D0 U33 ( .A1(inp[1]), .A2(rst_n), .Z(N48) );
  AN2D0 U34 ( .A1(inp[2]), .A2(rst_n), .Z(N49) );
  AN2D0 U35 ( .A1(inp[3]), .A2(rst_n), .Z(N50) );
  AN2D0 U36 ( .A1(inp[4]), .A2(rst_n), .Z(N51) );
  AN2D0 U37 ( .A1(inp[5]), .A2(rst_n), .Z(N52) );
  AN2D0 U38 ( .A1(inp[6]), .A2(rst_n), .Z(N53) );
  AN2D0 U39 ( .A1(inp[7]), .A2(rst_n), .Z(N54) );
  AN2D0 U40 ( .A1(inp[8]), .A2(rst_n), .Z(N55) );
  AN2D0 U41 ( .A1(inp[9]), .A2(rst_n), .Z(N56) );
  AN2D0 U42 ( .A1(inp[10]), .A2(rst_n), .Z(N57) );
  AN2D0 U43 ( .A1(inp[11]), .A2(rst_n), .Z(N58) );
  AN2D0 U44 ( .A1(inp[12]), .A2(rst_n), .Z(N59) );
  AN2D0 U45 ( .A1(inp[13]), .A2(rst_n), .Z(N60) );
  AN2D0 U46 ( .A1(inp[14]), .A2(rst_n), .Z(N61) );
  AN2D0 U47 ( .A1(inp[15]), .A2(rst_n), .Z(N62) );
  ND2D1 U48 ( .A1(n41), .A2(n42), .ZN(N68) );
  AOI22D0 U49 ( .A1(\mem2[1][0] ), .A2(n1), .B1(\mem2[4][0] ), .B2(n2), .ZN(
        n41) );
  AOI222D0 U50 ( .A1(\mem2[2][0] ), .A2(n3), .B1(\mem2[0][0] ), .B2(n4), .C1(
        \mem2[3][0] ), .C2(n5), .ZN(n42) );
  ND2D1 U51 ( .A1(n39), .A2(n40), .ZN(N69) );
  AOI22D0 U52 ( .A1(\mem2[1][1] ), .A2(n1), .B1(\mem2[4][1] ), .B2(n2), .ZN(
        n39) );
  AOI222D0 U53 ( .A1(\mem2[2][1] ), .A2(n3), .B1(\mem2[0][1] ), .B2(n4), .C1(
        \mem2[3][1] ), .C2(n5), .ZN(n40) );
  ND2D1 U54 ( .A1(n37), .A2(n38), .ZN(N70) );
  AOI22D0 U55 ( .A1(\mem2[1][2] ), .A2(n1), .B1(\mem2[4][2] ), .B2(n2), .ZN(
        n37) );
  AOI222D0 U56 ( .A1(\mem2[2][2] ), .A2(n3), .B1(\mem2[0][2] ), .B2(n4), .C1(
        \mem2[3][2] ), .C2(n5), .ZN(n38) );
  ND2D1 U57 ( .A1(n35), .A2(n36), .ZN(N71) );
  AOI22D0 U58 ( .A1(\mem2[1][3] ), .A2(n1), .B1(\mem2[4][3] ), .B2(n2), .ZN(
        n35) );
  AOI222D0 U59 ( .A1(\mem2[2][3] ), .A2(n3), .B1(\mem2[0][3] ), .B2(n4), .C1(
        \mem2[3][3] ), .C2(n5), .ZN(n36) );
  ND2D1 U60 ( .A1(n33), .A2(n34), .ZN(N72) );
  AOI22D0 U61 ( .A1(\mem2[1][4] ), .A2(n1), .B1(\mem2[4][4] ), .B2(n2), .ZN(
        n33) );
  AOI222D0 U62 ( .A1(\mem2[2][4] ), .A2(n3), .B1(\mem2[0][4] ), .B2(n4), .C1(
        \mem2[3][4] ), .C2(n5), .ZN(n34) );
  ND2D1 U63 ( .A1(n31), .A2(n32), .ZN(N73) );
  AOI22D0 U64 ( .A1(\mem2[1][5] ), .A2(n1), .B1(\mem2[4][5] ), .B2(n2), .ZN(
        n31) );
  AOI222D0 U65 ( .A1(\mem2[2][5] ), .A2(n3), .B1(\mem2[0][5] ), .B2(n4), .C1(
        \mem2[3][5] ), .C2(n5), .ZN(n32) );
  ND2D1 U66 ( .A1(n29), .A2(n30), .ZN(N74) );
  AOI22D0 U67 ( .A1(\mem2[1][6] ), .A2(n1), .B1(\mem2[4][6] ), .B2(n2), .ZN(
        n29) );
  AOI222D0 U68 ( .A1(\mem2[2][6] ), .A2(n3), .B1(\mem2[0][6] ), .B2(n4), .C1(
        \mem2[3][6] ), .C2(n5), .ZN(n30) );
  ND2D1 U69 ( .A1(n27), .A2(n28), .ZN(N75) );
  AOI22D0 U70 ( .A1(\mem2[1][7] ), .A2(n1), .B1(\mem2[4][7] ), .B2(n2), .ZN(
        n27) );
  AOI222D0 U71 ( .A1(\mem2[2][7] ), .A2(n3), .B1(\mem2[0][7] ), .B2(n4), .C1(
        \mem2[3][7] ), .C2(n5), .ZN(n28) );
  ND2D1 U72 ( .A1(n25), .A2(n26), .ZN(N76) );
  AOI22D0 U73 ( .A1(\mem2[1][8] ), .A2(n1), .B1(\mem2[4][8] ), .B2(n2), .ZN(
        n25) );
  AOI222D0 U74 ( .A1(\mem2[2][8] ), .A2(n3), .B1(\mem2[0][8] ), .B2(n4), .C1(
        \mem2[3][8] ), .C2(n5), .ZN(n26) );
  ND2D1 U75 ( .A1(n23), .A2(n24), .ZN(N77) );
  AOI22D0 U76 ( .A1(\mem2[1][9] ), .A2(n1), .B1(\mem2[4][9] ), .B2(n2), .ZN(
        n23) );
  AOI222D0 U77 ( .A1(\mem2[2][9] ), .A2(n3), .B1(\mem2[0][9] ), .B2(n4), .C1(
        \mem2[3][9] ), .C2(n5), .ZN(n24) );
  ND2D1 U78 ( .A1(n21), .A2(n22), .ZN(N78) );
  AOI22D0 U79 ( .A1(\mem2[1][10] ), .A2(n1), .B1(\mem2[4][10] ), .B2(n2), .ZN(
        n21) );
  AOI222D0 U80 ( .A1(\mem2[2][10] ), .A2(n3), .B1(\mem2[0][10] ), .B2(n4), 
        .C1(\mem2[3][10] ), .C2(n5), .ZN(n22) );
  ND2D1 U81 ( .A1(n19), .A2(n20), .ZN(N79) );
  AOI22D0 U82 ( .A1(\mem2[1][11] ), .A2(n1), .B1(\mem2[4][11] ), .B2(n2), .ZN(
        n19) );
  AOI222D0 U83 ( .A1(\mem2[2][11] ), .A2(n3), .B1(\mem2[0][11] ), .B2(n4), 
        .C1(\mem2[3][11] ), .C2(n5), .ZN(n20) );
  ND2D1 U84 ( .A1(n17), .A2(n18), .ZN(N80) );
  AOI22D0 U85 ( .A1(\mem2[1][12] ), .A2(n1), .B1(\mem2[4][12] ), .B2(n2), .ZN(
        n17) );
  AOI222D0 U86 ( .A1(\mem2[2][12] ), .A2(n3), .B1(\mem2[0][12] ), .B2(n4), 
        .C1(\mem2[3][12] ), .C2(n5), .ZN(n18) );
  ND2D1 U87 ( .A1(n15), .A2(n16), .ZN(N81) );
  AOI22D0 U88 ( .A1(\mem2[1][13] ), .A2(n1), .B1(\mem2[4][13] ), .B2(n2), .ZN(
        n15) );
  AOI222D0 U89 ( .A1(\mem2[2][13] ), .A2(n3), .B1(\mem2[0][13] ), .B2(n4), 
        .C1(\mem2[3][13] ), .C2(n5), .ZN(n16) );
  ND2D1 U90 ( .A1(n13), .A2(n14), .ZN(N82) );
  AOI22D0 U91 ( .A1(\mem2[1][14] ), .A2(n1), .B1(\mem2[4][14] ), .B2(n2), .ZN(
        n13) );
  AOI222D0 U92 ( .A1(\mem2[2][14] ), .A2(n3), .B1(\mem2[0][14] ), .B2(n4), 
        .C1(\mem2[3][14] ), .C2(n5), .ZN(n14) );
  ND2D1 U93 ( .A1(n6), .A2(n7), .ZN(N83) );
  AOI22D0 U94 ( .A1(\mem2[1][15] ), .A2(n1), .B1(\mem2[4][15] ), .B2(n2), .ZN(
        n6) );
  AOI222D0 U95 ( .A1(\mem2[2][15] ), .A2(n3), .B1(\mem2[0][15] ), .B2(n4), 
        .C1(\mem2[3][15] ), .C2(n5), .ZN(n7) );
endmodule


module Delayline_CB_DW01_inc_0 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;

  wire   [31:2] carry;

  CMPE22D1 U1_1_30 ( .A(A[30]), .B(carry[30]), .CO(carry[31]), .S(SUM[30]) );
  CMPE22D1 U1_1_27 ( .A(A[27]), .B(carry[27]), .CO(carry[28]), .S(SUM[27]) );
  CMPE22D1 U1_1_23 ( .A(A[23]), .B(carry[23]), .CO(carry[24]), .S(SUM[23]) );
  CMPE22D1 U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  CMPE22D1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  CMPE22D1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  CMPE22D1 U1_1_29 ( .A(A[29]), .B(carry[29]), .CO(carry[30]), .S(SUM[29]) );
  CMPE22D1 U1_1_26 ( .A(A[26]), .B(carry[26]), .CO(carry[27]), .S(SUM[26]) );
  CMPE22D1 U1_1_25 ( .A(A[25]), .B(carry[25]), .CO(carry[26]), .S(SUM[25]) );
  CMPE22D1 U1_1_22 ( .A(A[22]), .B(carry[22]), .CO(carry[23]), .S(SUM[22]) );
  CMPE22D1 U1_1_21 ( .A(A[21]), .B(carry[21]), .CO(carry[22]), .S(SUM[21]) );
  CMPE22D1 U1_1_19 ( .A(A[19]), .B(carry[19]), .CO(carry[20]), .S(SUM[19]) );
  CMPE22D1 U1_1_18 ( .A(A[18]), .B(carry[18]), .CO(carry[19]), .S(SUM[18]) );
  CMPE22D1 U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  CMPE22D1 U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  CMPE22D1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  CMPE22D1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  CMPE22D1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  CMPE22D1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  CMPE22D1 U1_1_28 ( .A(A[28]), .B(carry[28]), .CO(carry[29]), .S(SUM[28]) );
  CMPE22D1 U1_1_24 ( .A(A[24]), .B(carry[24]), .CO(carry[25]), .S(SUM[24]) );
  CMPE22D1 U1_1_20 ( .A(A[20]), .B(carry[20]), .CO(carry[21]), .S(SUM[20]) );
  CMPE22D1 U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  CMPE22D1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  CMPE22D1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  CMPE22D1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  CMPE22D1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  CMPE22D1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  CMPE22D1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  CMPE22D1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INVD1 U1 ( .I(A[0]), .ZN(SUM[0]) );
  CKXOR2D0 U2 ( .A1(carry[31]), .A2(A[31]), .Z(SUM[31]) );
endmodule


module Delayline_CB_DW01_dec_0 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  INVD1 U1 ( .I(A[12]), .ZN(n4) );
  INVD1 U2 ( .I(A[8]), .ZN(n2) );
  INVD1 U3 ( .I(A[10]), .ZN(n3) );
  INVD1 U4 ( .I(A[27]), .ZN(n5) );
  INVD1 U5 ( .I(A[29]), .ZN(n6) );
  INVD1 U6 ( .I(A[0]), .ZN(SUM[0]) );
  AO21D0 U7 ( .A1(n7), .A2(A[9]), .B(n8), .Z(SUM[9]) );
  OAI21D0 U8 ( .A1(n9), .A2(n2), .B(n7), .ZN(SUM[8]) );
  AO21D0 U9 ( .A1(n10), .A2(A[7]), .B(n9), .Z(SUM[7]) );
  IOA21D0 U10 ( .A1(n11), .A2(A[6]), .B(n10), .ZN(SUM[6]) );
  IOA21D0 U11 ( .A1(n12), .A2(A[5]), .B(n11), .ZN(SUM[5]) );
  IOA21D0 U12 ( .A1(n13), .A2(A[4]), .B(n12), .ZN(SUM[4]) );
  IOA21D0 U13 ( .A1(n14), .A2(A[3]), .B(n13), .ZN(SUM[3]) );
  CKXOR2D0 U14 ( .A1(A[31]), .A2(n15), .Z(SUM[31]) );
  NR2D0 U15 ( .A1(A[30]), .A2(n16), .ZN(n15) );
  XNR2D0 U16 ( .A1(n16), .A2(A[30]), .ZN(SUM[30]) );
  IOA21D0 U17 ( .A1(n17), .A2(A[2]), .B(n14), .ZN(SUM[2]) );
  OAI21D0 U18 ( .A1(n18), .A2(n6), .B(n16), .ZN(SUM[29]) );
  ND2D0 U19 ( .A1(n18), .A2(n6), .ZN(n16) );
  AO21D0 U20 ( .A1(n19), .A2(A[28]), .B(n18), .Z(SUM[28]) );
  NR2D0 U21 ( .A1(n19), .A2(A[28]), .ZN(n18) );
  OAI21D0 U22 ( .A1(n20), .A2(n5), .B(n19), .ZN(SUM[27]) );
  ND2D0 U23 ( .A1(n20), .A2(n5), .ZN(n19) );
  AO21D0 U24 ( .A1(n21), .A2(A[26]), .B(n20), .Z(SUM[26]) );
  NR2D0 U25 ( .A1(n21), .A2(A[26]), .ZN(n20) );
  IOA21D0 U26 ( .A1(n22), .A2(A[25]), .B(n21), .ZN(SUM[25]) );
  OR2D0 U27 ( .A1(n22), .A2(A[25]), .Z(n21) );
  IOA21D0 U28 ( .A1(n23), .A2(A[24]), .B(n22), .ZN(SUM[24]) );
  OR2D0 U29 ( .A1(n23), .A2(A[24]), .Z(n22) );
  IOA21D0 U30 ( .A1(n24), .A2(A[23]), .B(n23), .ZN(SUM[23]) );
  OR2D0 U31 ( .A1(n24), .A2(A[23]), .Z(n23) );
  IOA21D0 U32 ( .A1(n25), .A2(A[22]), .B(n24), .ZN(SUM[22]) );
  OR2D0 U33 ( .A1(n25), .A2(A[22]), .Z(n24) );
  IOA21D0 U34 ( .A1(n26), .A2(A[21]), .B(n25), .ZN(SUM[21]) );
  OR2D0 U35 ( .A1(n26), .A2(A[21]), .Z(n25) );
  IOA21D0 U36 ( .A1(n27), .A2(A[20]), .B(n26), .ZN(SUM[20]) );
  OR2D0 U37 ( .A1(n27), .A2(A[20]), .Z(n26) );
  IOA21D0 U38 ( .A1(A[0]), .A2(A[1]), .B(n17), .ZN(SUM[1]) );
  IOA21D0 U39 ( .A1(n28), .A2(A[19]), .B(n27), .ZN(SUM[19]) );
  OR2D0 U40 ( .A1(n28), .A2(A[19]), .Z(n27) );
  IOA21D0 U41 ( .A1(n29), .A2(A[18]), .B(n28), .ZN(SUM[18]) );
  OR2D0 U42 ( .A1(n29), .A2(A[18]), .Z(n28) );
  IOA21D0 U43 ( .A1(n30), .A2(A[17]), .B(n29), .ZN(SUM[17]) );
  OR2D0 U44 ( .A1(n30), .A2(A[17]), .Z(n29) );
  IOA21D0 U45 ( .A1(n31), .A2(A[16]), .B(n30), .ZN(SUM[16]) );
  OR2D0 U46 ( .A1(n31), .A2(A[16]), .Z(n30) );
  IOA21D0 U47 ( .A1(n32), .A2(A[15]), .B(n31), .ZN(SUM[15]) );
  OR2D0 U48 ( .A1(n32), .A2(A[15]), .Z(n31) );
  IOA21D0 U49 ( .A1(n33), .A2(A[14]), .B(n32), .ZN(SUM[14]) );
  OR2D0 U50 ( .A1(n33), .A2(A[14]), .Z(n32) );
  IOA21D0 U51 ( .A1(n34), .A2(A[13]), .B(n33), .ZN(SUM[13]) );
  OR2D0 U52 ( .A1(n34), .A2(A[13]), .Z(n33) );
  OAI21D0 U53 ( .A1(n35), .A2(n4), .B(n34), .ZN(SUM[12]) );
  ND2D0 U54 ( .A1(n35), .A2(n4), .ZN(n34) );
  AO21D0 U55 ( .A1(n36), .A2(A[11]), .B(n35), .Z(SUM[11]) );
  NR2D0 U56 ( .A1(n36), .A2(A[11]), .ZN(n35) );
  OAI21D0 U57 ( .A1(n8), .A2(n3), .B(n36), .ZN(SUM[10]) );
  ND2D0 U58 ( .A1(n8), .A2(n3), .ZN(n36) );
  NR2D0 U59 ( .A1(n7), .A2(A[9]), .ZN(n8) );
  ND2D0 U60 ( .A1(n9), .A2(n2), .ZN(n7) );
  NR2D0 U61 ( .A1(n10), .A2(A[7]), .ZN(n9) );
  OR2D0 U62 ( .A1(n11), .A2(A[6]), .Z(n10) );
  OR2D0 U63 ( .A1(n12), .A2(A[5]), .Z(n11) );
  OR2D0 U64 ( .A1(n13), .A2(A[4]), .Z(n12) );
  OR2D0 U65 ( .A1(n14), .A2(A[3]), .Z(n13) );
  OR2D0 U66 ( .A1(n17), .A2(A[2]), .Z(n14) );
  OR2D0 U67 ( .A1(A[1]), .A2(A[0]), .Z(n17) );
endmodule


module Delayline_CB ( rst_n, clk, sample_clk, sample, sample_out );
  input [15:0] sample;
  output [15:0] sample_out;
  input rst_n, clk, sample_clk;
  wire   rws_wire, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20,
         N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34,
         N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48,
         N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62,
         N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N74, N75, N76, N77,
         N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91,
         N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104,
         N105, N138, N139, N140, N141, N142, N143, N144, N145, N146, N147,
         N148, N149, N150, N151, N152, N153, N154, N155, N156, N157, N158,
         N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169,
         N170, N171, N172, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n1, n2, n24, n25, n26,
         n27, n28;
  wire   [2:0] adrs_wire;
  wire   [15:0] sample_write;
  wire   [31:0] counter;
  wire   [31:0] pointer;

  OR4D1 U37 ( .A1(pointer[24]), .A2(pointer[25]), .A3(pointer[26]), .A4(
        pointer[27]), .Z(n8) );
  OR4D1 U38 ( .A1(pointer[28]), .A2(pointer[29]), .A3(pointer[2]), .A4(
        pointer[30]), .Z(n7) );
  OR4D1 U39 ( .A1(pointer[31]), .A2(pointer[3]), .A3(pointer[4]), .A4(
        pointer[5]), .Z(n6) );
  OR4D1 U40 ( .A1(pointer[6]), .A2(pointer[7]), .A3(pointer[8]), .A4(
        pointer[9]), .Z(n5) );
  OR4D1 U42 ( .A1(pointer[0]), .A2(pointer[10]), .A3(pointer[11]), .A4(
        pointer[12]), .Z(n12) );
  OR4D1 U43 ( .A1(pointer[13]), .A2(pointer[14]), .A3(pointer[15]), .A4(
        pointer[16]), .Z(n11) );
  OR4D1 U44 ( .A1(pointer[17]), .A2(pointer[18]), .A3(pointer[19]), .A4(
        pointer[1]), .Z(n10) );
  OR4D1 U45 ( .A1(pointer[20]), .A2(pointer[21]), .A3(pointer[22]), .A4(
        pointer[23]), .Z(n9) );
  IAO21D1 U81 ( .A1(n14), .A2(n15), .B(n25), .ZN(n13) );
  SRAM U30_CBRAM ( .rst_n(rst_n), .rws(rws_wire), .addrs(adrs_wire), .inp(
        sample_write), .outp(sample_out) );
  Delayline_CB_DW01_inc_0 add_78 ( .A(counter), .SUM({N105, N104, N103, N102, 
        N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, 
        N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74})
         );
  Delayline_CB_DW01_dec_0 sub_67 ( .A(pointer), .SUM({N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, 
        N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9}) );
  EDFCNQD1 \sample_write_reg[15]  ( .D(sample[15]), .E(n25), .CP(clk), .CDN(
        rst_n), .Q(sample_write[15]) );
  EDFCNQD1 \sample_write_reg[14]  ( .D(sample[14]), .E(n25), .CP(clk), .CDN(
        rst_n), .Q(sample_write[14]) );
  EDFCNQD1 \sample_write_reg[13]  ( .D(sample[13]), .E(n25), .CP(clk), .CDN(
        rst_n), .Q(sample_write[13]) );
  EDFCNQD1 \sample_write_reg[12]  ( .D(sample[12]), .E(n25), .CP(clk), .CDN(
        rst_n), .Q(sample_write[12]) );
  EDFCNQD1 \sample_write_reg[11]  ( .D(sample[11]), .E(n25), .CP(clk), .CDN(
        rst_n), .Q(sample_write[11]) );
  EDFCNQD1 \sample_write_reg[10]  ( .D(sample[10]), .E(n25), .CP(clk), .CDN(
        rst_n), .Q(sample_write[10]) );
  EDFCNQD1 \sample_write_reg[9]  ( .D(sample[9]), .E(n25), .CP(clk), .CDN(
        rst_n), .Q(sample_write[9]) );
  EDFCNQD1 \sample_write_reg[8]  ( .D(sample[8]), .E(n25), .CP(clk), .CDN(
        rst_n), .Q(sample_write[8]) );
  EDFCNQD1 \sample_write_reg[7]  ( .D(sample[7]), .E(n25), .CP(clk), .CDN(
        rst_n), .Q(sample_write[7]) );
  EDFCNQD1 \sample_write_reg[6]  ( .D(sample[6]), .E(n25), .CP(clk), .CDN(
        rst_n), .Q(sample_write[6]) );
  EDFCNQD1 \sample_write_reg[5]  ( .D(sample[5]), .E(n25), .CP(clk), .CDN(
        rst_n), .Q(sample_write[5]) );
  EDFCNQD1 \sample_write_reg[4]  ( .D(sample[4]), .E(n25), .CP(clk), .CDN(
        rst_n), .Q(sample_write[4]) );
  EDFCNQD1 \sample_write_reg[3]  ( .D(sample[3]), .E(n25), .CP(clk), .CDN(
        rst_n), .Q(sample_write[3]) );
  EDFCNQD1 \sample_write_reg[2]  ( .D(sample[2]), .E(n25), .CP(clk), .CDN(
        rst_n), .Q(sample_write[2]) );
  EDFCNQD1 \sample_write_reg[1]  ( .D(sample[1]), .E(n25), .CP(clk), .CDN(
        rst_n), .Q(sample_write[1]) );
  EDFCNQD1 \sample_write_reg[0]  ( .D(sample[0]), .E(n25), .CP(clk), .CDN(
        rst_n), .Q(sample_write[0]) );
  DFSND1 rws_wire_reg ( .D(n26), .CP(clk), .SDN(rst_n), .Q(rws_wire) );
  DFCNQD1 \adrs_wire_reg[2]  ( .D(N172), .CP(clk), .CDN(rst_n), .Q(
        adrs_wire[2]) );
  DFCNQD1 \adrs_wire_reg[1]  ( .D(N171), .CP(clk), .CDN(rst_n), .Q(
        adrs_wire[1]) );
  DFCNQD1 \adrs_wire_reg[0]  ( .D(N170), .CP(clk), .CDN(rst_n), .Q(
        adrs_wire[0]) );
  DFCNQD1 \counter_reg[31]  ( .D(N169), .CP(clk), .CDN(rst_n), .Q(counter[31])
         );
  DFCNQD1 \counter_reg[23]  ( .D(N161), .CP(clk), .CDN(rst_n), .Q(counter[23])
         );
  DFCNQD1 \counter_reg[27]  ( .D(N165), .CP(clk), .CDN(rst_n), .Q(counter[27])
         );
  DFCNQD1 \counter_reg[19]  ( .D(N157), .CP(clk), .CDN(rst_n), .Q(counter[19])
         );
  DFCNQD1 \counter_reg[22]  ( .D(N160), .CP(clk), .CDN(rst_n), .Q(counter[22])
         );
  DFCNQD1 \counter_reg[26]  ( .D(N164), .CP(clk), .CDN(rst_n), .Q(counter[26])
         );
  DFCNQD1 \counter_reg[30]  ( .D(N168), .CP(clk), .CDN(rst_n), .Q(counter[30])
         );
  DFCNQD1 \counter_reg[18]  ( .D(N156), .CP(clk), .CDN(rst_n), .Q(counter[18])
         );
  DFCNQD1 \counter_reg[21]  ( .D(N159), .CP(clk), .CDN(rst_n), .Q(counter[21])
         );
  DFCNQD1 \counter_reg[25]  ( .D(N163), .CP(clk), .CDN(rst_n), .Q(counter[25])
         );
  DFCNQD1 \counter_reg[29]  ( .D(N167), .CP(clk), .CDN(rst_n), .Q(counter[29])
         );
  DFCNQD1 \counter_reg[20]  ( .D(N158), .CP(clk), .CDN(rst_n), .Q(counter[20])
         );
  DFCNQD1 \counter_reg[24]  ( .D(N162), .CP(clk), .CDN(rst_n), .Q(counter[24])
         );
  DFCNQD1 \counter_reg[28]  ( .D(N166), .CP(clk), .CDN(rst_n), .Q(counter[28])
         );
  DFCNQD1 \counter_reg[6]  ( .D(N144), .CP(clk), .CDN(rst_n), .Q(counter[6])
         );
  DFCNQD1 \counter_reg[12]  ( .D(N150), .CP(clk), .CDN(rst_n), .Q(counter[12])
         );
  DFCNQD1 \counter_reg[16]  ( .D(N154), .CP(clk), .CDN(rst_n), .Q(counter[16])
         );
  DFCNQD1 \counter_reg[5]  ( .D(N143), .CP(clk), .CDN(rst_n), .Q(counter[5])
         );
  DFCNQD1 \counter_reg[9]  ( .D(N147), .CP(clk), .CDN(rst_n), .Q(counter[9])
         );
  DFCNQD1 \counter_reg[15]  ( .D(N153), .CP(clk), .CDN(rst_n), .Q(counter[15])
         );
  DFCNQD1 \counter_reg[4]  ( .D(N142), .CP(clk), .CDN(rst_n), .Q(counter[4])
         );
  DFCNQD1 \counter_reg[8]  ( .D(N146), .CP(clk), .CDN(rst_n), .Q(counter[8])
         );
  DFCNQD1 \counter_reg[14]  ( .D(N152), .CP(clk), .CDN(rst_n), .Q(counter[14])
         );
  DFCNQD1 \counter_reg[3]  ( .D(N141), .CP(clk), .CDN(rst_n), .Q(counter[3])
         );
  DFCNQD1 \counter_reg[7]  ( .D(N145), .CP(clk), .CDN(rst_n), .Q(counter[7])
         );
  DFCNQD1 \counter_reg[13]  ( .D(N151), .CP(clk), .CDN(rst_n), .Q(counter[13])
         );
  DFCNQD1 \counter_reg[17]  ( .D(N155), .CP(clk), .CDN(rst_n), .Q(counter[17])
         );
  DFCNQD1 \counter_reg[10]  ( .D(N148), .CP(clk), .CDN(rst_n), .Q(counter[10])
         );
  DFCNQD1 \counter_reg[11]  ( .D(N149), .CP(clk), .CDN(rst_n), .Q(counter[11])
         );
  DFCNQD1 \counter_reg[2]  ( .D(N140), .CP(clk), .CDN(rst_n), .Q(counter[2])
         );
  DFCNQD1 \counter_reg[1]  ( .D(N139), .CP(clk), .CDN(rst_n), .Q(counter[1])
         );
  DFCNQD1 \counter_reg[0]  ( .D(N138), .CP(clk), .CDN(rst_n), .Q(counter[0])
         );
  EDFCNQD1 \pointer_reg[2]  ( .D(N43), .E(sample_clk), .CP(clk), .CDN(rst_n), 
        .Q(pointer[2]) );
  EDFCNQD1 \pointer_reg[4]  ( .D(N45), .E(sample_clk), .CP(clk), .CDN(rst_n), 
        .Q(pointer[4]) );
  EDFCNQD1 \pointer_reg[3]  ( .D(N44), .E(sample_clk), .CP(clk), .CDN(rst_n), 
        .Q(pointer[3]) );
  EDFCNQD1 \pointer_reg[1]  ( .D(N42), .E(sample_clk), .CP(clk), .CDN(rst_n), 
        .Q(pointer[1]) );
  EDFCNQD1 \pointer_reg[0]  ( .D(N41), .E(sample_clk), .CP(clk), .CDN(rst_n), 
        .Q(pointer[0]) );
  EDFCNQD1 \pointer_reg[5]  ( .D(N46), .E(sample_clk), .CP(clk), .CDN(rst_n), 
        .Q(pointer[5]) );
  EDFCNQD1 \pointer_reg[6]  ( .D(N47), .E(sample_clk), .CP(clk), .CDN(rst_n), 
        .Q(pointer[6]) );
  EDFCNQD1 \pointer_reg[7]  ( .D(N48), .E(sample_clk), .CP(clk), .CDN(rst_n), 
        .Q(pointer[7]) );
  EDFCNQD1 \pointer_reg[8]  ( .D(N49), .E(sample_clk), .CP(clk), .CDN(rst_n), 
        .Q(pointer[8]) );
  EDFCNQD1 \pointer_reg[9]  ( .D(N50), .E(sample_clk), .CP(clk), .CDN(rst_n), 
        .Q(pointer[9]) );
  EDFCNQD1 \pointer_reg[10]  ( .D(N51), .E(sample_clk), .CP(clk), .CDN(rst_n), 
        .Q(pointer[10]) );
  EDFCNQD1 \pointer_reg[11]  ( .D(N52), .E(sample_clk), .CP(clk), .CDN(rst_n), 
        .Q(pointer[11]) );
  EDFCNQD1 \pointer_reg[12]  ( .D(N53), .E(sample_clk), .CP(clk), .CDN(rst_n), 
        .Q(pointer[12]) );
  EDFCNQD1 \pointer_reg[13]  ( .D(N54), .E(sample_clk), .CP(clk), .CDN(rst_n), 
        .Q(pointer[13]) );
  EDFCNQD1 \pointer_reg[14]  ( .D(N55), .E(sample_clk), .CP(clk), .CDN(rst_n), 
        .Q(pointer[14]) );
  EDFCNQD1 \pointer_reg[15]  ( .D(N56), .E(sample_clk), .CP(clk), .CDN(rst_n), 
        .Q(pointer[15]) );
  EDFCNQD1 \pointer_reg[16]  ( .D(N57), .E(sample_clk), .CP(clk), .CDN(rst_n), 
        .Q(pointer[16]) );
  EDFCNQD1 \pointer_reg[17]  ( .D(N58), .E(sample_clk), .CP(clk), .CDN(rst_n), 
        .Q(pointer[17]) );
  EDFCNQD1 \pointer_reg[18]  ( .D(N59), .E(sample_clk), .CP(clk), .CDN(rst_n), 
        .Q(pointer[18]) );
  EDFCNQD1 \pointer_reg[19]  ( .D(N60), .E(sample_clk), .CP(clk), .CDN(rst_n), 
        .Q(pointer[19]) );
  EDFCNQD1 \pointer_reg[20]  ( .D(N61), .E(sample_clk), .CP(clk), .CDN(rst_n), 
        .Q(pointer[20]) );
  EDFCNQD1 \pointer_reg[21]  ( .D(N62), .E(sample_clk), .CP(clk), .CDN(rst_n), 
        .Q(pointer[21]) );
  EDFCNQD1 \pointer_reg[22]  ( .D(N63), .E(sample_clk), .CP(clk), .CDN(rst_n), 
        .Q(pointer[22]) );
  EDFCNQD1 \pointer_reg[23]  ( .D(N64), .E(sample_clk), .CP(clk), .CDN(rst_n), 
        .Q(pointer[23]) );
  EDFCNQD1 \pointer_reg[24]  ( .D(N65), .E(sample_clk), .CP(clk), .CDN(rst_n), 
        .Q(pointer[24]) );
  EDFCNQD1 \pointer_reg[25]  ( .D(N66), .E(sample_clk), .CP(clk), .CDN(rst_n), 
        .Q(pointer[25]) );
  EDFCNQD1 \pointer_reg[26]  ( .D(N67), .E(sample_clk), .CP(clk), .CDN(rst_n), 
        .Q(pointer[26]) );
  EDFCNQD1 \pointer_reg[27]  ( .D(N68), .E(sample_clk), .CP(clk), .CDN(rst_n), 
        .Q(pointer[27]) );
  EDFCNQD1 \pointer_reg[28]  ( .D(N69), .E(sample_clk), .CP(clk), .CDN(rst_n), 
        .Q(pointer[28]) );
  EDFCNQD1 \pointer_reg[29]  ( .D(N70), .E(sample_clk), .CP(clk), .CDN(rst_n), 
        .Q(pointer[29]) );
  EDFCNQD1 \pointer_reg[30]  ( .D(N71), .E(sample_clk), .CP(clk), .CDN(rst_n), 
        .Q(pointer[30]) );
  EDFCNQD1 \pointer_reg[31]  ( .D(N72), .E(sample_clk), .CP(clk), .CDN(rst_n), 
        .Q(pointer[31]) );
  ND2D1 U3 ( .A1(n3), .A2(n4), .ZN(n1) );
  BUFFD0 U4 ( .I(n27), .Z(n26) );
  INVD1 U5 ( .I(n13), .ZN(n24) );
  INVD1 U6 ( .I(n26), .ZN(n25) );
  INVD1 U7 ( .I(n24), .ZN(n2) );
  AN2D0 U8 ( .A1(N38), .A2(n1), .Z(N70) );
  AN2D0 U9 ( .A1(N36), .A2(n1), .Z(N68) );
  AN2D0 U10 ( .A1(N21), .A2(n1), .Z(N53) );
  AN2D0 U11 ( .A1(N19), .A2(n1), .Z(N51) );
  AN2D0 U12 ( .A1(N17), .A2(n1), .Z(N49) );
  ND4D1 U13 ( .A1(n20), .A2(n21), .A3(n22), .A4(n23), .ZN(n14) );
  ND4D1 U14 ( .A1(n16), .A2(n17), .A3(n18), .A4(n19), .ZN(n15) );
  NR4D0 U15 ( .A1(n5), .A2(n6), .A3(n7), .A4(n8), .ZN(n4) );
  NR4D0 U16 ( .A1(n9), .A2(n10), .A3(n11), .A4(n12), .ZN(n3) );
  BUFFD0 U17 ( .I(n28), .Z(n27) );
  AN2D0 U18 ( .A1(N37), .A2(n1), .Z(N69) );
  AN2D0 U19 ( .A1(N40), .A2(n1), .Z(N72) );
  AN2D0 U20 ( .A1(N39), .A2(n1), .Z(N71) );
  AN2D0 U21 ( .A1(N35), .A2(n1), .Z(N67) );
  AN2D0 U22 ( .A1(N34), .A2(n1), .Z(N66) );
  AN2D0 U23 ( .A1(N33), .A2(n1), .Z(N65) );
  AN2D0 U24 ( .A1(N32), .A2(n1), .Z(N64) );
  AN2D0 U25 ( .A1(N31), .A2(n1), .Z(N63) );
  AN2D0 U26 ( .A1(N30), .A2(n1), .Z(N62) );
  AN2D0 U27 ( .A1(N29), .A2(n1), .Z(N61) );
  AN2D0 U28 ( .A1(N28), .A2(n1), .Z(N60) );
  AN2D0 U29 ( .A1(N27), .A2(n1), .Z(N59) );
  AN2D0 U30 ( .A1(N26), .A2(n1), .Z(N58) );
  AO22D0 U31 ( .A1(sample_clk), .A2(pointer[31]), .B1(N105), .B2(n13), .Z(N169) );
  AO22D0 U32 ( .A1(sample_clk), .A2(pointer[30]), .B1(N104), .B2(n13), .Z(N168) );
  AO22D0 U33 ( .A1(sample_clk), .A2(pointer[29]), .B1(N103), .B2(n2), .Z(N167)
         );
  AO22D0 U34 ( .A1(sample_clk), .A2(pointer[28]), .B1(N102), .B2(n13), .Z(N166) );
  AO22D0 U35 ( .A1(sample_clk), .A2(pointer[27]), .B1(N101), .B2(n2), .Z(N165)
         );
  AO22D0 U36 ( .A1(sample_clk), .A2(pointer[26]), .B1(N100), .B2(n13), .Z(N164) );
  AO22D0 U41 ( .A1(sample_clk), .A2(pointer[25]), .B1(N99), .B2(n13), .Z(N163)
         );
  AO22D0 U46 ( .A1(sample_clk), .A2(pointer[24]), .B1(N98), .B2(n13), .Z(N162)
         );
  AO22D0 U47 ( .A1(sample_clk), .A2(pointer[23]), .B1(N97), .B2(n13), .Z(N161)
         );
  AO22D0 U48 ( .A1(sample_clk), .A2(pointer[22]), .B1(N96), .B2(n13), .Z(N160)
         );
  AO22D0 U49 ( .A1(sample_clk), .A2(pointer[21]), .B1(N95), .B2(n2), .Z(N159)
         );
  AO22D0 U50 ( .A1(sample_clk), .A2(pointer[20]), .B1(N94), .B2(n2), .Z(N158)
         );
  AO22D0 U51 ( .A1(n25), .A2(pointer[19]), .B1(N93), .B2(n2), .Z(N157) );
  AO22D0 U52 ( .A1(n25), .A2(pointer[18]), .B1(N92), .B2(n2), .Z(N156) );
  AO22D0 U53 ( .A1(sample_clk), .A2(pointer[17]), .B1(N91), .B2(n2), .Z(N155)
         );
  AO22D0 U54 ( .A1(n25), .A2(pointer[16]), .B1(N90), .B2(n2), .Z(N154) );
  AO22D0 U55 ( .A1(n25), .A2(pointer[15]), .B1(N89), .B2(n2), .Z(N153) );
  AN2D0 U56 ( .A1(N25), .A2(n1), .Z(N57) );
  AN2D0 U57 ( .A1(N24), .A2(n1), .Z(N56) );
  AN2D0 U58 ( .A1(N23), .A2(n1), .Z(N55) );
  AN2D0 U59 ( .A1(N22), .A2(n1), .Z(N54) );
  AN2D0 U60 ( .A1(N20), .A2(n1), .Z(N52) );
  AN2D0 U61 ( .A1(N18), .A2(n1), .Z(N50) );
  AN2D0 U62 ( .A1(N16), .A2(n1), .Z(N48) );
  NR4D0 U63 ( .A1(counter[26]), .A2(counter[25]), .A3(counter[24]), .A4(
        counter[23]), .ZN(n20) );
  NR4D0 U64 ( .A1(counter[22]), .A2(counter[21]), .A3(counter[20]), .A4(
        counter[1]), .ZN(n19) );
  NR4D0 U65 ( .A1(counter[19]), .A2(counter[18]), .A3(counter[17]), .A4(
        counter[16]), .ZN(n18) );
  NR4D0 U66 ( .A1(counter[9]), .A2(counter[8]), .A3(counter[7]), .A4(
        counter[6]), .ZN(n23) );
  NR4D0 U67 ( .A1(counter[5]), .A2(counter[4]), .A3(counter[3]), .A4(
        counter[31]), .ZN(n22) );
  NR4D0 U68 ( .A1(counter[15]), .A2(counter[14]), .A3(counter[13]), .A4(
        counter[12]), .ZN(n17) );
  NR4D0 U69 ( .A1(counter[30]), .A2(counter[29]), .A3(counter[28]), .A4(
        counter[27]), .ZN(n21) );
  INR4D0 U70 ( .A1(counter[2]), .B1(counter[11]), .B2(counter[10]), .B3(
        counter[0]), .ZN(n16) );
  AN2D0 U71 ( .A1(N15), .A2(n1), .Z(N47) );
  AO22D0 U72 ( .A1(sample_clk), .A2(pointer[0]), .B1(n26), .B2(counter[0]), 
        .Z(N170) );
  AO22D0 U73 ( .A1(n25), .A2(pointer[1]), .B1(n26), .B2(counter[1]), .Z(N171)
         );
  AO22D0 U74 ( .A1(n25), .A2(pointer[2]), .B1(n26), .B2(counter[2]), .Z(N172)
         );
  AO22D0 U75 ( .A1(sample_clk), .A2(pointer[14]), .B1(N88), .B2(n2), .Z(N152)
         );
  AO22D0 U76 ( .A1(n25), .A2(pointer[13]), .B1(N87), .B2(n2), .Z(N151) );
  AO22D0 U77 ( .A1(n25), .A2(pointer[12]), .B1(N86), .B2(n2), .Z(N150) );
  AO22D0 U78 ( .A1(sample_clk), .A2(pointer[11]), .B1(N85), .B2(n2), .Z(N149)
         );
  AO22D0 U79 ( .A1(n25), .A2(pointer[10]), .B1(N84), .B2(n2), .Z(N148) );
  AO22D0 U80 ( .A1(n25), .A2(pointer[9]), .B1(N83), .B2(n13), .Z(N147) );
  AO22D0 U82 ( .A1(sample_clk), .A2(pointer[8]), .B1(N82), .B2(n13), .Z(N146)
         );
  AO22D0 U83 ( .A1(n25), .A2(pointer[7]), .B1(N81), .B2(n13), .Z(N145) );
  AO22D0 U84 ( .A1(n25), .A2(pointer[6]), .B1(N80), .B2(n13), .Z(N144) );
  AO22D0 U85 ( .A1(n25), .A2(pointer[5]), .B1(N79), .B2(n13), .Z(N143) );
  AO22D0 U86 ( .A1(n25), .A2(pointer[4]), .B1(N78), .B2(n13), .Z(N142) );
  AO22D0 U87 ( .A1(sample_clk), .A2(pointer[3]), .B1(N77), .B2(n13), .Z(N141)
         );
  AO22D0 U88 ( .A1(n25), .A2(pointer[2]), .B1(N76), .B2(n13), .Z(N140) );
  AO22D0 U89 ( .A1(sample_clk), .A2(pointer[1]), .B1(N75), .B2(n13), .Z(N139)
         );
  AO22D0 U90 ( .A1(n25), .A2(pointer[0]), .B1(N74), .B2(n13), .Z(N138) );
  IND2D1 U91 ( .A1(N11), .B1(n1), .ZN(N43) );
  AN2D0 U92 ( .A1(N9), .A2(n1), .Z(N41) );
  AN2D0 U93 ( .A1(N14), .A2(n1), .Z(N46) );
  AN2D0 U94 ( .A1(N13), .A2(n1), .Z(N45) );
  AN2D0 U95 ( .A1(N12), .A2(n1), .Z(N44) );
  AN2D0 U96 ( .A1(N10), .A2(n1), .Z(N42) );
  INVD1 U97 ( .I(sample_clk), .ZN(n28) );
endmodule


module FIR_Processor_DW01_dec_0 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  INVD1 U1 ( .I(A[10]), .ZN(n3) );
  INVD1 U2 ( .I(A[8]), .ZN(n2) );
  INVD1 U3 ( .I(A[12]), .ZN(n4) );
  INVD1 U4 ( .I(A[29]), .ZN(n6) );
  INVD1 U5 ( .I(A[27]), .ZN(n5) );
  INVD1 U6 ( .I(A[0]), .ZN(SUM[0]) );
  AO21D0 U7 ( .A1(n7), .A2(A[9]), .B(n8), .Z(SUM[9]) );
  OAI21D0 U8 ( .A1(n9), .A2(n2), .B(n7), .ZN(SUM[8]) );
  AO21D0 U9 ( .A1(n10), .A2(A[7]), .B(n9), .Z(SUM[7]) );
  IOA21D0 U10 ( .A1(n11), .A2(A[6]), .B(n10), .ZN(SUM[6]) );
  IOA21D0 U11 ( .A1(n12), .A2(A[5]), .B(n11), .ZN(SUM[5]) );
  IOA21D0 U12 ( .A1(n13), .A2(A[4]), .B(n12), .ZN(SUM[4]) );
  IOA21D0 U13 ( .A1(n14), .A2(A[3]), .B(n13), .ZN(SUM[3]) );
  CKXOR2D0 U14 ( .A1(A[31]), .A2(n15), .Z(SUM[31]) );
  NR2D0 U15 ( .A1(A[30]), .A2(n16), .ZN(n15) );
  XNR2D0 U16 ( .A1(n16), .A2(A[30]), .ZN(SUM[30]) );
  IOA21D0 U17 ( .A1(n17), .A2(A[2]), .B(n14), .ZN(SUM[2]) );
  OAI21D0 U18 ( .A1(n18), .A2(n6), .B(n16), .ZN(SUM[29]) );
  ND2D0 U19 ( .A1(n18), .A2(n6), .ZN(n16) );
  AO21D0 U20 ( .A1(n19), .A2(A[28]), .B(n18), .Z(SUM[28]) );
  NR2D0 U21 ( .A1(n19), .A2(A[28]), .ZN(n18) );
  OAI21D0 U22 ( .A1(n20), .A2(n5), .B(n19), .ZN(SUM[27]) );
  ND2D0 U23 ( .A1(n20), .A2(n5), .ZN(n19) );
  AO21D0 U24 ( .A1(n21), .A2(A[26]), .B(n20), .Z(SUM[26]) );
  NR2D0 U25 ( .A1(n21), .A2(A[26]), .ZN(n20) );
  IOA21D0 U26 ( .A1(n22), .A2(A[25]), .B(n21), .ZN(SUM[25]) );
  OR2D0 U27 ( .A1(n22), .A2(A[25]), .Z(n21) );
  IOA21D0 U28 ( .A1(n23), .A2(A[24]), .B(n22), .ZN(SUM[24]) );
  OR2D0 U29 ( .A1(n23), .A2(A[24]), .Z(n22) );
  IOA21D0 U30 ( .A1(n24), .A2(A[23]), .B(n23), .ZN(SUM[23]) );
  OR2D0 U31 ( .A1(n24), .A2(A[23]), .Z(n23) );
  IOA21D0 U32 ( .A1(n25), .A2(A[22]), .B(n24), .ZN(SUM[22]) );
  OR2D0 U33 ( .A1(n25), .A2(A[22]), .Z(n24) );
  IOA21D0 U34 ( .A1(n26), .A2(A[21]), .B(n25), .ZN(SUM[21]) );
  OR2D0 U35 ( .A1(n26), .A2(A[21]), .Z(n25) );
  IOA21D0 U36 ( .A1(n27), .A2(A[20]), .B(n26), .ZN(SUM[20]) );
  OR2D0 U37 ( .A1(n27), .A2(A[20]), .Z(n26) );
  IOA21D0 U38 ( .A1(A[0]), .A2(A[1]), .B(n17), .ZN(SUM[1]) );
  IOA21D0 U39 ( .A1(n28), .A2(A[19]), .B(n27), .ZN(SUM[19]) );
  OR2D0 U40 ( .A1(n28), .A2(A[19]), .Z(n27) );
  IOA21D0 U41 ( .A1(n29), .A2(A[18]), .B(n28), .ZN(SUM[18]) );
  OR2D0 U42 ( .A1(n29), .A2(A[18]), .Z(n28) );
  IOA21D0 U43 ( .A1(n30), .A2(A[17]), .B(n29), .ZN(SUM[17]) );
  OR2D0 U44 ( .A1(n30), .A2(A[17]), .Z(n29) );
  IOA21D0 U45 ( .A1(n31), .A2(A[16]), .B(n30), .ZN(SUM[16]) );
  OR2D0 U46 ( .A1(n31), .A2(A[16]), .Z(n30) );
  IOA21D0 U47 ( .A1(n32), .A2(A[15]), .B(n31), .ZN(SUM[15]) );
  OR2D0 U48 ( .A1(n32), .A2(A[15]), .Z(n31) );
  IOA21D0 U49 ( .A1(n33), .A2(A[14]), .B(n32), .ZN(SUM[14]) );
  OR2D0 U50 ( .A1(n33), .A2(A[14]), .Z(n32) );
  IOA21D0 U51 ( .A1(n34), .A2(A[13]), .B(n33), .ZN(SUM[13]) );
  OR2D0 U52 ( .A1(n34), .A2(A[13]), .Z(n33) );
  OAI21D0 U53 ( .A1(n35), .A2(n4), .B(n34), .ZN(SUM[12]) );
  ND2D0 U54 ( .A1(n35), .A2(n4), .ZN(n34) );
  AO21D0 U55 ( .A1(n36), .A2(A[11]), .B(n35), .Z(SUM[11]) );
  NR2D0 U56 ( .A1(n36), .A2(A[11]), .ZN(n35) );
  OAI21D0 U57 ( .A1(n8), .A2(n3), .B(n36), .ZN(SUM[10]) );
  ND2D0 U58 ( .A1(n8), .A2(n3), .ZN(n36) );
  NR2D0 U59 ( .A1(n7), .A2(A[9]), .ZN(n8) );
  ND2D0 U60 ( .A1(n9), .A2(n2), .ZN(n7) );
  NR2D0 U61 ( .A1(n10), .A2(A[7]), .ZN(n9) );
  OR2D0 U62 ( .A1(n11), .A2(A[6]), .Z(n10) );
  OR2D0 U63 ( .A1(n12), .A2(A[5]), .Z(n11) );
  OR2D0 U64 ( .A1(n13), .A2(A[4]), .Z(n12) );
  OR2D0 U65 ( .A1(n14), .A2(A[3]), .Z(n13) );
  OR2D0 U66 ( .A1(n17), .A2(A[2]), .Z(n14) );
  OR2D0 U67 ( .A1(A[1]), .A2(A[0]), .Z(n17) );
endmodule


module FIR_Processor_DW_mult_uns_0 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n83, n84, n86, n87, n88, n89, n90, n91, n92, n93, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n295, n296, n297, n298, n299, n300, n301, n302,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904;

  CMPE32D1 U53 ( .A(n84), .B(n88), .CI(n53), .CO(n52), .S(product[30]) );
  CMPE32D1 U54 ( .A(n89), .B(n91), .CI(n54), .CO(n53), .S(product[29]) );
  CMPE32D1 U55 ( .A(n92), .B(n96), .CI(n55), .CO(n54), .S(product[28]) );
  CMPE32D1 U56 ( .A(n97), .B(n101), .CI(n56), .CO(n55), .S(product[27]) );
  CMPE32D1 U57 ( .A(n102), .B(n108), .CI(n57), .CO(n56), .S(product[26]) );
  CMPE32D1 U58 ( .A(n109), .B(n114), .CI(n58), .CO(n57), .S(product[25]) );
  CMPE32D1 U59 ( .A(n115), .B(n122), .CI(n59), .CO(n58), .S(product[24]) );
  CMPE32D1 U60 ( .A(n123), .B(n130), .CI(n60), .CO(n59), .S(product[23]) );
  CMPE32D1 U61 ( .A(n131), .B(n140), .CI(n61), .CO(n60), .S(product[22]) );
  CMPE32D1 U62 ( .A(n141), .B(n149), .CI(n62), .CO(n61), .S(product[21]) );
  CMPE32D1 U63 ( .A(n150), .B(n160), .CI(n63), .CO(n62), .S(product[20]) );
  CMPE32D1 U64 ( .A(n161), .B(n171), .CI(n64), .CO(n63), .S(product[19]) );
  CMPE32D1 U65 ( .A(n172), .B(n184), .CI(n65), .CO(n64), .S(product[18]) );
  CMPE32D1 U66 ( .A(n185), .B(n196), .CI(n66), .CO(n65), .S(product[17]) );
  CMPE32D1 U67 ( .A(n197), .B(n207), .CI(n67), .CO(n66), .S(product[16]) );
  CMPE32D1 U68 ( .A(n218), .B(n208), .CI(n68), .CO(n67), .S(product[15]) );
  CMPE32D1 U69 ( .A(n227), .B(n219), .CI(n69), .CO(n68), .S(product[14]) );
  CMPE32D1 U70 ( .A(n228), .B(n237), .CI(n70), .CO(n69), .S(product[13]) );
  CMPE32D1 U71 ( .A(n245), .B(n238), .CI(n71), .CO(n70), .S(product[12]) );
  CMPE32D1 U72 ( .A(n253), .B(n246), .CI(n72), .CO(n71), .S(product[11]) );
  CMPE32D1 U73 ( .A(n259), .B(n254), .CI(n73), .CO(n72), .S(product[10]) );
  CMPE32D1 U74 ( .A(n266), .B(n260), .CI(n74), .CO(n73), .S(product[9]) );
  CMPE32D1 U75 ( .A(n271), .B(n267), .CI(n75), .CO(n74), .S(product[8]) );
  CMPE32D1 U76 ( .A(n276), .B(n272), .CI(n76), .CO(n75), .S(product[7]) );
  CMPE32D1 U77 ( .A(n278), .B(n277), .CI(n77), .CO(n76), .S(product[6]) );
  CMPE32D1 U78 ( .A(n282), .B(n279), .CI(n78), .CO(n77), .S(product[5]) );
  CMPE32D1 U79 ( .A(n284), .B(n283), .CI(n79), .CO(n78), .S(product[4]) );
  CMPE32D1 U80 ( .A(n292), .B(n285), .CI(n80), .CO(n79), .S(product[3]) );
  CMPE32D1 U81 ( .A(n428), .B(n444), .CI(n81), .CO(n80), .S(product[2]) );
  CMPE22D1 U82 ( .A(n293), .B(n445), .CO(n81), .S(product[1]) );
  CMPE32D1 U84 ( .A(n86), .B(n304), .CI(n87), .CO(n83), .S(n84) );
  CMPE42D1 U86 ( .A(n93), .B(n295), .C(n321), .CIX(n90), .D(n305), .CO(n88), 
        .COX(n87), .S(n89) );
  CMPE42D1 U87 ( .A(n734), .B(n322), .C(n306), .CIX(n95), .D(n98), .CO(n91), 
        .COX(n90), .S(n92) );
  CMPE42D1 U89 ( .A(n323), .B(n307), .C(n99), .CIX(n100), .D(n103), .CO(n96), 
        .COX(n95), .S(n97) );
  CMPE32D1 U90 ( .A(n105), .B(n296), .CI(n339), .CO(n98), .S(n99) );
  CMPE42D1 U91 ( .A(n308), .B(n110), .C(n104), .CIX(n107), .D(n111), .CO(n101), 
        .COX(n100), .S(n102) );
  CMPE32D1 U92 ( .A(n729), .B(n324), .CI(n340), .CO(n103), .S(n104) );
  CMPE42D1 U94 ( .A(n341), .B(n116), .C(n112), .CIX(n113), .D(n117), .CO(n108), 
        .COX(n107), .S(n109) );
  CMPE42D1 U95 ( .A(n119), .B(n297), .C(n357), .CIX(n309), .D(n325), .CO(n111), 
        .COX(n110), .S(n112) );
  CMPE42D1 U96 ( .A(n310), .B(n124), .C(n118), .CIX(n121), .D(n125), .CO(n114), 
        .COX(n113), .S(n115) );
  CMPE42D1 U97 ( .A(n730), .B(n358), .C(n342), .CIX(n127), .D(n326), .CO(n117), 
        .COX(n116), .S(n118) );
  CMPE42D1 U99 ( .A(n311), .B(n135), .C(n126), .CIX(n129), .D(n133), .CO(n122), 
        .COX(n121), .S(n123) );
  CMPE42D1 U100 ( .A(n327), .B(n359), .C(n343), .CIX(n132), .D(n128), .CO(n125), .COX(n124), .S(n126) );
  CMPE32D1 U101 ( .A(n137), .B(n298), .CI(n375), .CO(n127), .S(n128) );
  CMPE42D1 U102 ( .A(n136), .B(n146), .C(n134), .CIX(n139), .D(n143), .CO(n130), .COX(n129), .S(n131) );
  CMPE42D1 U103 ( .A(n312), .B(n360), .C(n344), .CIX(n142), .D(n145), .CO(n133), .COX(n132), .S(n134) );
  CMPE32D1 U104 ( .A(n731), .B(n376), .CI(n328), .CO(n135), .S(n136) );
  CMPE42D1 U106 ( .A(n147), .B(n155), .C(n152), .CIX(n148), .D(n144), .CO(n140), .COX(n139), .S(n141) );
  CMPE42D1 U107 ( .A(n361), .B(n329), .C(n345), .CIX(n151), .D(n154), .CO(n143), .COX(n142), .S(n144) );
  CMPE42D1 U108 ( .A(n157), .B(n299), .C(n393), .CIX(n313), .D(n377), .CO(n146), .COX(n145), .S(n147) );
  CMPE42D1 U109 ( .A(n156), .B(n166), .C(n163), .CIX(n159), .D(n153), .CO(n149), .COX(n148), .S(n150) );
  CMPE42D1 U110 ( .A(n362), .B(n330), .C(n346), .CIX(n165), .D(n162), .CO(n152), .COX(n151), .S(n153) );
  CMPE42D1 U111 ( .A(n732), .B(n394), .C(n378), .CIX(n168), .D(n314), .CO(n155), .COX(n154), .S(n156) );
  CMPE42D1 U113 ( .A(n164), .B(n167), .C(n174), .CIX(n170), .D(n177), .CO(n160), .COX(n159), .S(n161) );
  CMPE42D1 U114 ( .A(n315), .B(n347), .C(n363), .CIX(n173), .D(n179), .CO(n163), .COX(n162), .S(n164) );
  CMPE42D1 U115 ( .A(n331), .B(n395), .C(n379), .CIX(n176), .D(n169), .CO(n166), .COX(n165), .S(n167) );
  CMPE32D1 U116 ( .A(n181), .B(n300), .CI(n411), .CO(n168), .S(n169) );
  CMPE42D1 U117 ( .A(n178), .B(n190), .C(n175), .CIX(n183), .D(n187), .CO(n171), .COX(n170), .S(n172) );
  CMPE42D1 U118 ( .A(n364), .B(n316), .C(n332), .CIX(n186), .D(n180), .CO(n174), .COX(n173), .S(n175) );
  CMPE42D1 U119 ( .A(n348), .B(n396), .C(n380), .CIX(n189), .D(n192), .CO(n177), .COX(n176), .S(n178) );
  CMPE32D1 U120 ( .A(n301), .B(n733), .CI(n412), .CO(n179), .S(n180) );
  CMPE42D1 U122 ( .A(n191), .B(n199), .C(n202), .CIX(n195), .D(n188), .CO(n184), .COX(n183), .S(n185) );
  CMPE42D1 U123 ( .A(n349), .B(n317), .C(n204), .CIX(n198), .D(n193), .CO(n187), .COX(n186), .S(n188) );
  CMPE42D1 U124 ( .A(n333), .B(n397), .C(n381), .CIX(n201), .D(n365), .CO(n190), .COX(n189), .S(n191) );
  CMPE32D1 U125 ( .A(n733), .B(n742), .CI(n413), .CO(n192), .S(n193) );
  CMPE42D1 U127 ( .A(n203), .B(n210), .C(n213), .CIX(n206), .D(n200), .CO(n196), .COX(n195), .S(n197) );
  CMPE42D1 U128 ( .A(n382), .B(n318), .C(n366), .CIX(n209), .D(n205), .CO(n199), .COX(n198), .S(n200) );
  CMPE42D1 U129 ( .A(n350), .B(n414), .C(n398), .CIX(n212), .D(n215), .CO(n202), .COX(n201), .S(n203) );
  CMPE32D1 U130 ( .A(n302), .B(n334), .CI(n430), .CO(n204), .S(n205) );
  CMPE42D1 U131 ( .A(n224), .B(n214), .C(n211), .CIX(n217), .D(n221), .CO(n207), .COX(n206), .S(n208) );
  CMPE42D1 U132 ( .A(n351), .B(n399), .C(n335), .CIX(n223), .D(n367), .CO(n210), .COX(n209), .S(n211) );
  CMPE42D1 U133 ( .A(n383), .B(n431), .C(n415), .CIX(n220), .D(n216), .CO(n213), .COX(n212), .S(n214) );
  CMPE22D1 U134 ( .A(n319), .B(n286), .CO(n215), .S(n216) );
  CMPE42D1 U135 ( .A(n232), .B(n225), .C(n222), .CIX(n226), .D(n230), .CO(n218), .COX(n217), .S(n219) );
  CMPE42D1 U136 ( .A(n416), .B(n368), .C(n400), .CIX(n229), .D(n384), .CO(n221), .COX(n220), .S(n222) );
  CMPE42D1 U137 ( .A(n320), .B(n352), .C(n432), .CIX(n234), .D(n336), .CO(n224), .COX(n223), .S(n225) );
  CMPE42D1 U138 ( .A(n242), .B(n233), .C(n231), .CIX(n236), .D(n240), .CO(n227), .COX(n226), .S(n228) );
  CMPE42D1 U139 ( .A(n417), .B(n369), .C(n401), .CIX(n239), .D(n235), .CO(n230), .COX(n229), .S(n231) );
  CMPE32D1 U140 ( .A(n385), .B(n433), .CI(n353), .CO(n232), .S(n233) );
  CMPE22D1 U141 ( .A(n337), .B(n287), .CO(n234), .S(n235) );
  CMPE42D1 U142 ( .A(n354), .B(n243), .C(n241), .CIX(n244), .D(n248), .CO(n237), .COX(n236), .S(n238) );
  CMPE42D1 U143 ( .A(n386), .B(n418), .C(n402), .CIX(n247), .D(n250), .CO(n240), .COX(n239), .S(n241) );
  CMPE32D1 U144 ( .A(n338), .B(n370), .CI(n434), .CO(n242), .S(n243) );
  CMPE42D1 U145 ( .A(n387), .B(n371), .C(n252), .CIX(n249), .D(n256), .CO(n245), .COX(n244), .S(n246) );
  CMPE42D1 U146 ( .A(n403), .B(n435), .C(n419), .CIX(n255), .D(n251), .CO(n248), .COX(n247), .S(n249) );
  CMPE22D1 U147 ( .A(n355), .B(n288), .CO(n250), .S(n251) );
  CMPE42D1 U148 ( .A(n420), .B(n404), .C(n261), .CIX(n257), .D(n258), .CO(n253), .COX(n252), .S(n254) );
  CMPE42D1 U149 ( .A(n356), .B(n388), .C(n436), .CIX(n263), .D(n372), .CO(n256), .COX(n255), .S(n257) );
  CMPE42D1 U150 ( .A(n437), .B(n264), .C(n268), .CIX(n265), .D(n262), .CO(n259), .COX(n258), .S(n260) );
  CMPE32D1 U151 ( .A(n405), .B(n389), .CI(n421), .CO(n261), .S(n262) );
  CMPE22D1 U152 ( .A(n373), .B(n289), .CO(n263), .S(n264) );
  CMPE42D1 U153 ( .A(n422), .B(n390), .C(n273), .CIX(n270), .D(n269), .CO(n266), .COX(n265), .S(n267) );
  CMPE32D1 U154 ( .A(n374), .B(n406), .CI(n438), .CO(n268), .S(n269) );
  CMPE42D1 U155 ( .A(n439), .B(n407), .C(n423), .CIX(n275), .D(n274), .CO(n271), .COX(n270), .S(n272) );
  CMPE22D1 U156 ( .A(n391), .B(n290), .CO(n273), .S(n274) );
  CMPE42D1 U157 ( .A(n392), .B(n440), .C(n424), .CIX(n280), .D(n408), .CO(n276), .COX(n275), .S(n277) );
  CMPE32D1 U158 ( .A(n441), .B(n425), .CI(n281), .CO(n278), .S(n279) );
  CMPE22D1 U159 ( .A(n409), .B(n291), .CO(n280), .S(n281) );
  CMPE32D1 U160 ( .A(n410), .B(n442), .CI(n426), .CO(n282), .S(n283) );
  CMPE22D1 U161 ( .A(n443), .B(n427), .CO(n284), .S(n285) );
  XNR2D1 U532 ( .A1(a[1]), .A2(a[2]), .ZN(n714) );
  XNR2D1 U533 ( .A1(a[3]), .A2(a[4]), .ZN(n715) );
  XNR2D1 U534 ( .A1(a[5]), .A2(a[6]), .ZN(n716) );
  XNR2D1 U535 ( .A1(a[7]), .A2(a[8]), .ZN(n717) );
  XNR2D1 U536 ( .A1(a[9]), .A2(a[10]), .ZN(n718) );
  XNR2D1 U537 ( .A1(a[11]), .A2(a[12]), .ZN(n719) );
  XNR2D1 U538 ( .A1(a[13]), .A2(a[14]), .ZN(n720) );
  BUFFD0 U539 ( .I(b[0]), .Z(n728) );
  INVD1 U540 ( .I(n181), .ZN(n733) );
  INVD1 U541 ( .I(b[2]), .ZN(n756) );
  INVD1 U542 ( .I(n157), .ZN(n732) );
  INVD1 U543 ( .I(b[1]), .ZN(n757) );
  INVD1 U544 ( .I(n728), .ZN(n758) );
  INVD1 U545 ( .I(n119), .ZN(n730) );
  INVD1 U546 ( .I(n93), .ZN(n734) );
  INVD1 U547 ( .I(n137), .ZN(n731) );
  INVD1 U548 ( .I(n105), .ZN(n729) );
  INVD1 U549 ( .I(b[3]), .ZN(n759) );
  INVD1 U550 ( .I(a[0]), .ZN(n743) );
  ND2D1 U551 ( .A1(a[1]), .A2(n743), .ZN(n764) );
  INVD1 U552 ( .I(a[3]), .ZN(n741) );
  INVD1 U553 ( .I(a[5]), .ZN(n740) );
  INVD1 U554 ( .I(a[7]), .ZN(n739) );
  INVD1 U555 ( .I(a[9]), .ZN(n738) );
  INVD1 U556 ( .I(a[11]), .ZN(n737) );
  INVD1 U557 ( .I(a[13]), .ZN(n736) );
  INVD1 U558 ( .I(a[1]), .ZN(n742) );
  INVD1 U559 ( .I(a[15]), .ZN(n735) );
  BUFFD0 U560 ( .I(n781), .Z(n721) );
  ND2D1 U561 ( .A1(n714), .A2(n898), .ZN(n781) );
  BUFFD0 U562 ( .I(n798), .Z(n722) );
  ND2D1 U563 ( .A1(n715), .A2(n899), .ZN(n798) );
  BUFFD0 U564 ( .I(n815), .Z(n723) );
  ND2D1 U565 ( .A1(n716), .A2(n900), .ZN(n815) );
  BUFFD0 U566 ( .I(n832), .Z(n724) );
  ND2D1 U567 ( .A1(n717), .A2(n901), .ZN(n832) );
  BUFFD0 U568 ( .I(n849), .Z(n725) );
  ND2D1 U569 ( .A1(n718), .A2(n902), .ZN(n849) );
  BUFFD0 U570 ( .I(n866), .Z(n726) );
  ND2D1 U571 ( .A1(n719), .A2(n903), .ZN(n866) );
  BUFFD0 U572 ( .I(n763), .Z(n727) );
  ND2D1 U573 ( .A1(n720), .A2(n904), .ZN(n763) );
  INVD1 U574 ( .I(b[4]), .ZN(n744) );
  INVD1 U575 ( .I(b[6]), .ZN(n746) );
  INVD1 U576 ( .I(b[8]), .ZN(n748) );
  INVD1 U577 ( .I(b[10]), .ZN(n750) );
  INVD1 U578 ( .I(b[12]), .ZN(n752) );
  INVD1 U579 ( .I(b[7]), .ZN(n747) );
  INVD1 U580 ( .I(b[11]), .ZN(n751) );
  INVD1 U581 ( .I(b[5]), .ZN(n745) );
  INVD1 U582 ( .I(b[9]), .ZN(n749) );
  INVD1 U583 ( .I(b[13]), .ZN(n753) );
  INVD1 U584 ( .I(b[15]), .ZN(n755) );
  INVD1 U585 ( .I(b[14]), .ZN(n754) );
  XNR3D0 U586 ( .A1(n760), .A2(n761), .A3(n762), .ZN(product[31]) );
  AOI21D0 U587 ( .A1(n727), .A2(n720), .B(n735), .ZN(n762) );
  XNR3D0 U588 ( .A1(n83), .A2(n52), .A3(n86), .ZN(n761) );
  NR2D0 U589 ( .A1(n735), .A2(n755), .ZN(n760) );
  NR2D0 U590 ( .A1(n743), .A2(n758), .ZN(product[0]) );
  NR2D0 U591 ( .A1(n752), .A2(n735), .ZN(n93) );
  ND2D0 U592 ( .A1(b[14]), .A2(a[15]), .ZN(n86) );
  OAI22D0 U593 ( .A1(n728), .A2(n764), .B1(n765), .B2(n743), .ZN(n445) );
  OAI22D0 U594 ( .A1(n765), .A2(n764), .B1(n766), .B2(n743), .ZN(n444) );
  XNR2D0 U595 ( .A1(n742), .A2(n757), .ZN(n765) );
  OAI22D0 U596 ( .A1(n766), .A2(n764), .B1(n767), .B2(n743), .ZN(n443) );
  XNR2D0 U597 ( .A1(n742), .A2(n756), .ZN(n766) );
  OAI22D0 U598 ( .A1(n767), .A2(n764), .B1(n768), .B2(n743), .ZN(n442) );
  XNR2D0 U599 ( .A1(n742), .A2(n759), .ZN(n767) );
  OAI22D0 U600 ( .A1(n768), .A2(n764), .B1(n769), .B2(n743), .ZN(n441) );
  XNR2D0 U601 ( .A1(n742), .A2(n744), .ZN(n768) );
  OAI22D0 U602 ( .A1(n769), .A2(n764), .B1(n770), .B2(n743), .ZN(n440) );
  XNR2D0 U603 ( .A1(n742), .A2(n745), .ZN(n769) );
  OAI22D0 U604 ( .A1(n770), .A2(n764), .B1(n771), .B2(n743), .ZN(n439) );
  XNR2D0 U605 ( .A1(n742), .A2(n746), .ZN(n770) );
  OAI22D0 U606 ( .A1(n771), .A2(n764), .B1(n772), .B2(n743), .ZN(n438) );
  XNR2D0 U607 ( .A1(n742), .A2(n747), .ZN(n771) );
  OAI22D0 U608 ( .A1(n772), .A2(n764), .B1(n773), .B2(n743), .ZN(n437) );
  XNR2D0 U609 ( .A1(n742), .A2(n748), .ZN(n772) );
  OAI22D0 U610 ( .A1(n773), .A2(n764), .B1(n774), .B2(n743), .ZN(n436) );
  XNR2D0 U611 ( .A1(n742), .A2(n749), .ZN(n773) );
  OAI22D0 U612 ( .A1(n774), .A2(n764), .B1(n775), .B2(n743), .ZN(n435) );
  XNR2D0 U613 ( .A1(n742), .A2(n750), .ZN(n774) );
  OAI22D0 U614 ( .A1(n775), .A2(n764), .B1(n776), .B2(n743), .ZN(n434) );
  XNR2D0 U615 ( .A1(n742), .A2(n751), .ZN(n775) );
  OAI22D0 U616 ( .A1(n776), .A2(n764), .B1(n777), .B2(n743), .ZN(n433) );
  XNR2D0 U617 ( .A1(n742), .A2(n752), .ZN(n776) );
  OAI22D0 U618 ( .A1(n777), .A2(n764), .B1(n778), .B2(n743), .ZN(n432) );
  XNR2D0 U619 ( .A1(n742), .A2(n753), .ZN(n777) );
  OAI22D0 U620 ( .A1(n778), .A2(n764), .B1(n779), .B2(n743), .ZN(n431) );
  XNR2D0 U621 ( .A1(n742), .A2(n754), .ZN(n778) );
  OAI22D0 U622 ( .A1(n779), .A2(n764), .B1(n742), .B2(n743), .ZN(n430) );
  XNR2D0 U623 ( .A1(n742), .A2(n755), .ZN(n779) );
  NR2D0 U624 ( .A1(n714), .A2(n758), .ZN(n428) );
  OAI22D0 U625 ( .A1(n780), .A2(n721), .B1(n714), .B2(n782), .ZN(n427) );
  XNR2D0 U626 ( .A1(n758), .A2(n741), .ZN(n780) );
  OAI22D0 U627 ( .A1(n782), .A2(n721), .B1(n714), .B2(n783), .ZN(n426) );
  XNR2D0 U628 ( .A1(n741), .A2(n757), .ZN(n782) );
  OAI22D0 U629 ( .A1(n783), .A2(n721), .B1(n714), .B2(n784), .ZN(n425) );
  XNR2D0 U630 ( .A1(n741), .A2(n756), .ZN(n783) );
  OAI22D0 U631 ( .A1(n784), .A2(n721), .B1(n714), .B2(n785), .ZN(n424) );
  XNR2D0 U632 ( .A1(n741), .A2(n759), .ZN(n784) );
  OAI22D0 U633 ( .A1(n785), .A2(n721), .B1(n714), .B2(n786), .ZN(n423) );
  XNR2D0 U634 ( .A1(n741), .A2(n744), .ZN(n785) );
  OAI22D0 U635 ( .A1(n786), .A2(n721), .B1(n714), .B2(n787), .ZN(n422) );
  XNR2D0 U636 ( .A1(n741), .A2(n745), .ZN(n786) );
  OAI22D0 U637 ( .A1(n787), .A2(n721), .B1(n714), .B2(n788), .ZN(n421) );
  XNR2D0 U638 ( .A1(n741), .A2(n746), .ZN(n787) );
  OAI22D0 U639 ( .A1(n788), .A2(n721), .B1(n714), .B2(n789), .ZN(n420) );
  XNR2D0 U640 ( .A1(n741), .A2(n747), .ZN(n788) );
  OAI22D0 U641 ( .A1(n789), .A2(n721), .B1(n714), .B2(n790), .ZN(n419) );
  XNR2D0 U642 ( .A1(n741), .A2(n748), .ZN(n789) );
  OAI22D0 U643 ( .A1(n790), .A2(n721), .B1(n714), .B2(n791), .ZN(n418) );
  XNR2D0 U644 ( .A1(n741), .A2(n749), .ZN(n790) );
  OAI22D0 U645 ( .A1(n791), .A2(n721), .B1(n714), .B2(n792), .ZN(n417) );
  XNR2D0 U646 ( .A1(n741), .A2(n750), .ZN(n791) );
  OAI22D0 U647 ( .A1(n792), .A2(n721), .B1(n714), .B2(n793), .ZN(n416) );
  XNR2D0 U648 ( .A1(n741), .A2(n751), .ZN(n792) );
  OAI22D0 U649 ( .A1(n793), .A2(n721), .B1(n714), .B2(n794), .ZN(n415) );
  XNR2D0 U650 ( .A1(n741), .A2(n752), .ZN(n793) );
  OAI22D0 U651 ( .A1(n794), .A2(n721), .B1(n714), .B2(n795), .ZN(n414) );
  XNR2D0 U652 ( .A1(n741), .A2(n753), .ZN(n794) );
  OAI22D0 U653 ( .A1(n795), .A2(n721), .B1(n714), .B2(n796), .ZN(n413) );
  XNR2D0 U654 ( .A1(n741), .A2(n754), .ZN(n795) );
  OAI22D0 U655 ( .A1(n796), .A2(n721), .B1(n714), .B2(n741), .ZN(n412) );
  XNR2D0 U656 ( .A1(n741), .A2(n755), .ZN(n796) );
  AO21D0 U657 ( .A1(n721), .A2(n714), .B(n741), .Z(n411) );
  NR2D0 U658 ( .A1(n715), .A2(n758), .ZN(n410) );
  OAI22D0 U659 ( .A1(n797), .A2(n722), .B1(n715), .B2(n799), .ZN(n409) );
  XNR2D0 U660 ( .A1(n758), .A2(n740), .ZN(n797) );
  OAI22D0 U661 ( .A1(n799), .A2(n722), .B1(n715), .B2(n800), .ZN(n408) );
  XNR2D0 U662 ( .A1(n740), .A2(n757), .ZN(n799) );
  OAI22D0 U663 ( .A1(n800), .A2(n722), .B1(n715), .B2(n801), .ZN(n407) );
  XNR2D0 U664 ( .A1(n740), .A2(n756), .ZN(n800) );
  OAI22D0 U665 ( .A1(n801), .A2(n722), .B1(n715), .B2(n802), .ZN(n406) );
  XNR2D0 U666 ( .A1(n740), .A2(n759), .ZN(n801) );
  OAI22D0 U667 ( .A1(n802), .A2(n722), .B1(n715), .B2(n803), .ZN(n405) );
  XNR2D0 U668 ( .A1(n740), .A2(n744), .ZN(n802) );
  OAI22D0 U669 ( .A1(n803), .A2(n722), .B1(n715), .B2(n804), .ZN(n404) );
  XNR2D0 U670 ( .A1(n740), .A2(n745), .ZN(n803) );
  OAI22D0 U671 ( .A1(n804), .A2(n722), .B1(n715), .B2(n805), .ZN(n403) );
  XNR2D0 U672 ( .A1(n740), .A2(n746), .ZN(n804) );
  OAI22D0 U673 ( .A1(n805), .A2(n722), .B1(n715), .B2(n806), .ZN(n402) );
  XNR2D0 U674 ( .A1(n740), .A2(n747), .ZN(n805) );
  OAI22D0 U675 ( .A1(n806), .A2(n722), .B1(n715), .B2(n807), .ZN(n401) );
  XNR2D0 U676 ( .A1(n740), .A2(n748), .ZN(n806) );
  OAI22D0 U677 ( .A1(n807), .A2(n722), .B1(n715), .B2(n808), .ZN(n400) );
  XNR2D0 U678 ( .A1(n740), .A2(n749), .ZN(n807) );
  OAI22D0 U679 ( .A1(n808), .A2(n722), .B1(n715), .B2(n809), .ZN(n399) );
  XNR2D0 U680 ( .A1(n740), .A2(n750), .ZN(n808) );
  OAI22D0 U681 ( .A1(n809), .A2(n722), .B1(n715), .B2(n810), .ZN(n398) );
  XNR2D0 U682 ( .A1(n740), .A2(n751), .ZN(n809) );
  OAI22D0 U683 ( .A1(n810), .A2(n722), .B1(n715), .B2(n811), .ZN(n397) );
  XNR2D0 U684 ( .A1(n740), .A2(n752), .ZN(n810) );
  OAI22D0 U685 ( .A1(n811), .A2(n722), .B1(n715), .B2(n812), .ZN(n396) );
  XNR2D0 U686 ( .A1(n740), .A2(n753), .ZN(n811) );
  OAI22D0 U687 ( .A1(n812), .A2(n722), .B1(n715), .B2(n813), .ZN(n395) );
  XNR2D0 U688 ( .A1(n740), .A2(n754), .ZN(n812) );
  OAI22D0 U689 ( .A1(n813), .A2(n722), .B1(n715), .B2(n740), .ZN(n394) );
  XNR2D0 U690 ( .A1(n740), .A2(n755), .ZN(n813) );
  AO21D0 U691 ( .A1(n722), .A2(n715), .B(n740), .Z(n393) );
  NR2D0 U692 ( .A1(n716), .A2(n758), .ZN(n392) );
  OAI22D0 U693 ( .A1(n814), .A2(n723), .B1(n716), .B2(n816), .ZN(n391) );
  XNR2D0 U694 ( .A1(n758), .A2(n739), .ZN(n814) );
  OAI22D0 U695 ( .A1(n816), .A2(n723), .B1(n716), .B2(n817), .ZN(n390) );
  XNR2D0 U696 ( .A1(n739), .A2(n757), .ZN(n816) );
  OAI22D0 U697 ( .A1(n817), .A2(n723), .B1(n716), .B2(n818), .ZN(n389) );
  XNR2D0 U698 ( .A1(n739), .A2(n756), .ZN(n817) );
  OAI22D0 U699 ( .A1(n818), .A2(n723), .B1(n716), .B2(n819), .ZN(n388) );
  XNR2D0 U700 ( .A1(n739), .A2(n759), .ZN(n818) );
  OAI22D0 U701 ( .A1(n819), .A2(n723), .B1(n716), .B2(n820), .ZN(n387) );
  XNR2D0 U702 ( .A1(n739), .A2(n744), .ZN(n819) );
  OAI22D0 U703 ( .A1(n820), .A2(n723), .B1(n716), .B2(n821), .ZN(n386) );
  XNR2D0 U704 ( .A1(n739), .A2(n745), .ZN(n820) );
  OAI22D0 U705 ( .A1(n821), .A2(n723), .B1(n716), .B2(n822), .ZN(n385) );
  XNR2D0 U706 ( .A1(n739), .A2(n746), .ZN(n821) );
  OAI22D0 U707 ( .A1(n822), .A2(n723), .B1(n716), .B2(n823), .ZN(n384) );
  XNR2D0 U708 ( .A1(n739), .A2(n747), .ZN(n822) );
  OAI22D0 U709 ( .A1(n823), .A2(n723), .B1(n716), .B2(n824), .ZN(n383) );
  XNR2D0 U710 ( .A1(n739), .A2(n748), .ZN(n823) );
  OAI22D0 U711 ( .A1(n824), .A2(n723), .B1(n716), .B2(n825), .ZN(n382) );
  XNR2D0 U712 ( .A1(n739), .A2(n749), .ZN(n824) );
  OAI22D0 U713 ( .A1(n825), .A2(n723), .B1(n716), .B2(n826), .ZN(n381) );
  XNR2D0 U714 ( .A1(n739), .A2(n750), .ZN(n825) );
  OAI22D0 U715 ( .A1(n826), .A2(n723), .B1(n716), .B2(n827), .ZN(n380) );
  XNR2D0 U716 ( .A1(n739), .A2(n751), .ZN(n826) );
  OAI22D0 U717 ( .A1(n827), .A2(n723), .B1(n716), .B2(n828), .ZN(n379) );
  XNR2D0 U718 ( .A1(n739), .A2(n752), .ZN(n827) );
  OAI22D0 U719 ( .A1(n828), .A2(n723), .B1(n716), .B2(n829), .ZN(n378) );
  XNR2D0 U720 ( .A1(n739), .A2(n753), .ZN(n828) );
  OAI22D0 U721 ( .A1(n829), .A2(n723), .B1(n716), .B2(n830), .ZN(n377) );
  XNR2D0 U722 ( .A1(n739), .A2(n754), .ZN(n829) );
  OAI22D0 U723 ( .A1(n830), .A2(n723), .B1(n716), .B2(n739), .ZN(n376) );
  XNR2D0 U724 ( .A1(n739), .A2(n755), .ZN(n830) );
  AO21D0 U725 ( .A1(n723), .A2(n716), .B(n739), .Z(n375) );
  NR2D0 U726 ( .A1(n717), .A2(n758), .ZN(n374) );
  OAI22D0 U727 ( .A1(n831), .A2(n724), .B1(n717), .B2(n833), .ZN(n373) );
  XNR2D0 U728 ( .A1(n758), .A2(n738), .ZN(n831) );
  OAI22D0 U729 ( .A1(n833), .A2(n724), .B1(n717), .B2(n834), .ZN(n372) );
  XNR2D0 U730 ( .A1(n738), .A2(n757), .ZN(n833) );
  OAI22D0 U731 ( .A1(n834), .A2(n724), .B1(n717), .B2(n835), .ZN(n371) );
  XNR2D0 U732 ( .A1(n738), .A2(n756), .ZN(n834) );
  OAI22D0 U733 ( .A1(n835), .A2(n724), .B1(n717), .B2(n836), .ZN(n370) );
  XNR2D0 U734 ( .A1(n738), .A2(n759), .ZN(n835) );
  OAI22D0 U735 ( .A1(n836), .A2(n724), .B1(n717), .B2(n837), .ZN(n369) );
  XNR2D0 U736 ( .A1(n738), .A2(n744), .ZN(n836) );
  OAI22D0 U737 ( .A1(n837), .A2(n724), .B1(n717), .B2(n838), .ZN(n368) );
  XNR2D0 U738 ( .A1(n738), .A2(n745), .ZN(n837) );
  OAI22D0 U739 ( .A1(n838), .A2(n724), .B1(n717), .B2(n839), .ZN(n367) );
  XNR2D0 U740 ( .A1(n738), .A2(n746), .ZN(n838) );
  OAI22D0 U741 ( .A1(n839), .A2(n724), .B1(n717), .B2(n840), .ZN(n366) );
  XNR2D0 U742 ( .A1(n738), .A2(n747), .ZN(n839) );
  OAI22D0 U743 ( .A1(n840), .A2(n724), .B1(n717), .B2(n841), .ZN(n365) );
  XNR2D0 U744 ( .A1(n738), .A2(n748), .ZN(n840) );
  OAI22D0 U745 ( .A1(n841), .A2(n724), .B1(n717), .B2(n842), .ZN(n364) );
  XNR2D0 U746 ( .A1(n738), .A2(n749), .ZN(n841) );
  OAI22D0 U747 ( .A1(n842), .A2(n724), .B1(n717), .B2(n843), .ZN(n363) );
  XNR2D0 U748 ( .A1(n738), .A2(n750), .ZN(n842) );
  OAI22D0 U749 ( .A1(n843), .A2(n724), .B1(n717), .B2(n844), .ZN(n362) );
  XNR2D0 U750 ( .A1(n738), .A2(n751), .ZN(n843) );
  OAI22D0 U751 ( .A1(n844), .A2(n724), .B1(n717), .B2(n845), .ZN(n361) );
  XNR2D0 U752 ( .A1(n738), .A2(n752), .ZN(n844) );
  OAI22D0 U753 ( .A1(n845), .A2(n724), .B1(n717), .B2(n846), .ZN(n360) );
  XNR2D0 U754 ( .A1(n738), .A2(n753), .ZN(n845) );
  OAI22D0 U755 ( .A1(n846), .A2(n724), .B1(n717), .B2(n847), .ZN(n359) );
  XNR2D0 U756 ( .A1(n738), .A2(n754), .ZN(n846) );
  OAI22D0 U757 ( .A1(n847), .A2(n724), .B1(n717), .B2(n738), .ZN(n358) );
  XNR2D0 U758 ( .A1(n738), .A2(n755), .ZN(n847) );
  AO21D0 U759 ( .A1(n724), .A2(n717), .B(n738), .Z(n357) );
  NR2D0 U760 ( .A1(n718), .A2(n758), .ZN(n356) );
  OAI22D0 U761 ( .A1(n848), .A2(n725), .B1(n718), .B2(n850), .ZN(n355) );
  XNR2D0 U762 ( .A1(n758), .A2(n737), .ZN(n848) );
  OAI22D0 U763 ( .A1(n850), .A2(n725), .B1(n718), .B2(n851), .ZN(n354) );
  XNR2D0 U764 ( .A1(n737), .A2(n757), .ZN(n850) );
  OAI22D0 U765 ( .A1(n851), .A2(n725), .B1(n718), .B2(n852), .ZN(n353) );
  XNR2D0 U766 ( .A1(n737), .A2(n756), .ZN(n851) );
  OAI22D0 U767 ( .A1(n852), .A2(n725), .B1(n718), .B2(n853), .ZN(n352) );
  XNR2D0 U768 ( .A1(n737), .A2(n759), .ZN(n852) );
  OAI22D0 U769 ( .A1(n853), .A2(n725), .B1(n718), .B2(n854), .ZN(n351) );
  XNR2D0 U770 ( .A1(n737), .A2(n744), .ZN(n853) );
  OAI22D0 U771 ( .A1(n854), .A2(n725), .B1(n718), .B2(n855), .ZN(n350) );
  XNR2D0 U772 ( .A1(n737), .A2(n745), .ZN(n854) );
  OAI22D0 U773 ( .A1(n855), .A2(n725), .B1(n718), .B2(n856), .ZN(n349) );
  XNR2D0 U774 ( .A1(n737), .A2(n746), .ZN(n855) );
  OAI22D0 U775 ( .A1(n856), .A2(n725), .B1(n718), .B2(n857), .ZN(n348) );
  XNR2D0 U776 ( .A1(n737), .A2(n747), .ZN(n856) );
  OAI22D0 U777 ( .A1(n857), .A2(n725), .B1(n718), .B2(n858), .ZN(n347) );
  XNR2D0 U778 ( .A1(n737), .A2(n748), .ZN(n857) );
  OAI22D0 U779 ( .A1(n858), .A2(n725), .B1(n718), .B2(n859), .ZN(n346) );
  XNR2D0 U780 ( .A1(n737), .A2(n749), .ZN(n858) );
  OAI22D0 U781 ( .A1(n859), .A2(n725), .B1(n718), .B2(n860), .ZN(n345) );
  XNR2D0 U782 ( .A1(n737), .A2(n750), .ZN(n859) );
  OAI22D0 U783 ( .A1(n860), .A2(n725), .B1(n718), .B2(n861), .ZN(n344) );
  XNR2D0 U784 ( .A1(n737), .A2(n751), .ZN(n860) );
  OAI22D0 U785 ( .A1(n861), .A2(n725), .B1(n718), .B2(n862), .ZN(n343) );
  XNR2D0 U786 ( .A1(n737), .A2(n752), .ZN(n861) );
  OAI22D0 U787 ( .A1(n862), .A2(n725), .B1(n718), .B2(n863), .ZN(n342) );
  XNR2D0 U788 ( .A1(n737), .A2(n753), .ZN(n862) );
  OAI22D0 U789 ( .A1(n863), .A2(n725), .B1(n718), .B2(n864), .ZN(n341) );
  XNR2D0 U790 ( .A1(n737), .A2(n754), .ZN(n863) );
  OAI22D0 U791 ( .A1(n864), .A2(n725), .B1(n718), .B2(n737), .ZN(n340) );
  XNR2D0 U792 ( .A1(n737), .A2(n755), .ZN(n864) );
  AO21D0 U793 ( .A1(n725), .A2(n718), .B(n737), .Z(n339) );
  NR2D0 U794 ( .A1(n719), .A2(n758), .ZN(n338) );
  OAI22D0 U795 ( .A1(n865), .A2(n726), .B1(n719), .B2(n867), .ZN(n337) );
  XNR2D0 U796 ( .A1(n758), .A2(n736), .ZN(n865) );
  OAI22D0 U797 ( .A1(n867), .A2(n726), .B1(n719), .B2(n868), .ZN(n336) );
  XNR2D0 U798 ( .A1(n736), .A2(n757), .ZN(n867) );
  OAI22D0 U799 ( .A1(n868), .A2(n726), .B1(n719), .B2(n869), .ZN(n335) );
  XNR2D0 U800 ( .A1(n736), .A2(n756), .ZN(n868) );
  OAI22D0 U801 ( .A1(n869), .A2(n726), .B1(n719), .B2(n870), .ZN(n334) );
  XNR2D0 U802 ( .A1(n736), .A2(n759), .ZN(n869) );
  OAI22D0 U803 ( .A1(n870), .A2(n726), .B1(n719), .B2(n871), .ZN(n333) );
  XNR2D0 U804 ( .A1(n736), .A2(n744), .ZN(n870) );
  OAI22D0 U805 ( .A1(n871), .A2(n726), .B1(n719), .B2(n872), .ZN(n332) );
  XNR2D0 U806 ( .A1(n736), .A2(n745), .ZN(n871) );
  OAI22D0 U807 ( .A1(n872), .A2(n726), .B1(n719), .B2(n873), .ZN(n331) );
  XNR2D0 U808 ( .A1(n736), .A2(n746), .ZN(n872) );
  OAI22D0 U809 ( .A1(n873), .A2(n726), .B1(n719), .B2(n874), .ZN(n330) );
  XNR2D0 U810 ( .A1(n736), .A2(n747), .ZN(n873) );
  OAI22D0 U811 ( .A1(n874), .A2(n726), .B1(n719), .B2(n875), .ZN(n329) );
  XNR2D0 U812 ( .A1(n736), .A2(n748), .ZN(n874) );
  OAI22D0 U813 ( .A1(n875), .A2(n726), .B1(n719), .B2(n876), .ZN(n328) );
  XNR2D0 U814 ( .A1(n736), .A2(n749), .ZN(n875) );
  OAI22D0 U815 ( .A1(n876), .A2(n726), .B1(n719), .B2(n877), .ZN(n327) );
  XNR2D0 U816 ( .A1(n736), .A2(n750), .ZN(n876) );
  OAI22D0 U817 ( .A1(n877), .A2(n726), .B1(n719), .B2(n878), .ZN(n326) );
  XNR2D0 U818 ( .A1(n736), .A2(n751), .ZN(n877) );
  OAI22D0 U819 ( .A1(n878), .A2(n726), .B1(n719), .B2(n879), .ZN(n325) );
  XNR2D0 U820 ( .A1(n736), .A2(n752), .ZN(n878) );
  OAI22D0 U821 ( .A1(n879), .A2(n726), .B1(n719), .B2(n880), .ZN(n324) );
  XNR2D0 U822 ( .A1(n736), .A2(n753), .ZN(n879) );
  OAI22D0 U823 ( .A1(n880), .A2(n726), .B1(n719), .B2(n881), .ZN(n323) );
  XNR2D0 U824 ( .A1(n736), .A2(n754), .ZN(n880) );
  OAI22D0 U825 ( .A1(n881), .A2(n726), .B1(n719), .B2(n736), .ZN(n322) );
  XNR2D0 U826 ( .A1(n736), .A2(n755), .ZN(n881) );
  AO21D0 U827 ( .A1(n726), .A2(n719), .B(n736), .Z(n321) );
  NR2D0 U828 ( .A1(n720), .A2(n758), .ZN(n320) );
  OAI22D0 U829 ( .A1(n882), .A2(n727), .B1(n720), .B2(n883), .ZN(n319) );
  XNR2D0 U830 ( .A1(n735), .A2(n758), .ZN(n882) );
  OAI22D0 U831 ( .A1(n883), .A2(n727), .B1(n720), .B2(n884), .ZN(n318) );
  XNR2D0 U832 ( .A1(n735), .A2(n757), .ZN(n883) );
  OAI22D0 U833 ( .A1(n884), .A2(n727), .B1(n720), .B2(n885), .ZN(n317) );
  XNR2D0 U834 ( .A1(n735), .A2(n756), .ZN(n884) );
  OAI22D0 U835 ( .A1(n885), .A2(n727), .B1(n720), .B2(n886), .ZN(n316) );
  XNR2D0 U836 ( .A1(n735), .A2(n759), .ZN(n885) );
  OAI22D0 U837 ( .A1(n886), .A2(n727), .B1(n720), .B2(n887), .ZN(n315) );
  XNR2D0 U838 ( .A1(n735), .A2(n744), .ZN(n886) );
  OAI22D0 U839 ( .A1(n887), .A2(n727), .B1(n720), .B2(n888), .ZN(n314) );
  XNR2D0 U840 ( .A1(n735), .A2(n745), .ZN(n887) );
  OAI22D0 U841 ( .A1(n888), .A2(n727), .B1(n720), .B2(n889), .ZN(n313) );
  XNR2D0 U842 ( .A1(n735), .A2(n746), .ZN(n888) );
  OAI22D0 U843 ( .A1(n889), .A2(n727), .B1(n720), .B2(n890), .ZN(n312) );
  XNR2D0 U844 ( .A1(n735), .A2(n747), .ZN(n889) );
  OAI22D0 U845 ( .A1(n890), .A2(n727), .B1(n720), .B2(n891), .ZN(n311) );
  XNR2D0 U846 ( .A1(n735), .A2(n748), .ZN(n890) );
  OAI22D0 U847 ( .A1(n891), .A2(n727), .B1(n720), .B2(n892), .ZN(n310) );
  XNR2D0 U848 ( .A1(n735), .A2(n749), .ZN(n891) );
  OAI22D0 U849 ( .A1(n892), .A2(n727), .B1(n720), .B2(n893), .ZN(n309) );
  XNR2D0 U850 ( .A1(n735), .A2(n750), .ZN(n892) );
  OAI22D0 U851 ( .A1(n893), .A2(n727), .B1(n720), .B2(n894), .ZN(n308) );
  XNR2D0 U852 ( .A1(n735), .A2(n751), .ZN(n893) );
  OAI22D0 U853 ( .A1(n894), .A2(n727), .B1(n720), .B2(n895), .ZN(n307) );
  XNR2D0 U854 ( .A1(n735), .A2(n752), .ZN(n894) );
  OAI22D0 U855 ( .A1(n895), .A2(n727), .B1(n720), .B2(n896), .ZN(n306) );
  XNR2D0 U856 ( .A1(n735), .A2(n753), .ZN(n895) );
  OAI22D0 U857 ( .A1(n896), .A2(n727), .B1(n720), .B2(n897), .ZN(n305) );
  XNR2D0 U858 ( .A1(n735), .A2(n754), .ZN(n896) );
  OAI22D0 U859 ( .A1(n897), .A2(n727), .B1(n720), .B2(n735), .ZN(n304) );
  XNR2D0 U860 ( .A1(n735), .A2(n755), .ZN(n897) );
  NR2D0 U861 ( .A1(n735), .A2(n758), .ZN(n302) );
  NR2D0 U862 ( .A1(n735), .A2(n756), .ZN(n301) );
  NR2D0 U863 ( .A1(n735), .A2(n759), .ZN(n300) );
  NR2D0 U864 ( .A1(n735), .A2(n745), .ZN(n299) );
  NR2D0 U865 ( .A1(n735), .A2(n747), .ZN(n298) );
  NR2D0 U866 ( .A1(n735), .A2(n749), .ZN(n297) );
  NR2D0 U867 ( .A1(n735), .A2(n751), .ZN(n296) );
  NR2D0 U868 ( .A1(n735), .A2(n753), .ZN(n295) );
  OAI21D0 U869 ( .A1(n728), .A2(n742), .B(n764), .ZN(n293) );
  OAI32D0 U870 ( .A1(n741), .A2(n728), .A3(n714), .B1(n741), .B2(n721), .ZN(
        n292) );
  XNR2D0 U871 ( .A1(n741), .A2(a[2]), .ZN(n898) );
  OAI32D0 U872 ( .A1(n740), .A2(n728), .A3(n715), .B1(n740), .B2(n722), .ZN(
        n291) );
  XNR2D0 U873 ( .A1(n740), .A2(a[4]), .ZN(n899) );
  OAI32D0 U874 ( .A1(n739), .A2(n728), .A3(n716), .B1(n739), .B2(n723), .ZN(
        n290) );
  XNR2D0 U875 ( .A1(n739), .A2(a[6]), .ZN(n900) );
  OAI32D0 U876 ( .A1(n738), .A2(n728), .A3(n717), .B1(n738), .B2(n724), .ZN(
        n289) );
  XNR2D0 U877 ( .A1(n738), .A2(a[8]), .ZN(n901) );
  OAI32D0 U878 ( .A1(n737), .A2(n728), .A3(n718), .B1(n737), .B2(n725), .ZN(
        n288) );
  XNR2D0 U879 ( .A1(n737), .A2(a[10]), .ZN(n902) );
  OAI32D0 U880 ( .A1(n736), .A2(n728), .A3(n719), .B1(n736), .B2(n726), .ZN(
        n287) );
  XNR2D0 U881 ( .A1(n736), .A2(a[12]), .ZN(n903) );
  OAI32D0 U882 ( .A1(n735), .A2(n728), .A3(n720), .B1(n735), .B2(n727), .ZN(
        n286) );
  XNR2D0 U883 ( .A1(n735), .A2(a[14]), .ZN(n904) );
  NR2D0 U884 ( .A1(n757), .A2(n735), .ZN(n181) );
  NR2D0 U885 ( .A1(n744), .A2(n735), .ZN(n157) );
  NR2D0 U886 ( .A1(n746), .A2(n735), .ZN(n137) );
  NR2D0 U887 ( .A1(n748), .A2(n735), .ZN(n119) );
  NR2D0 U888 ( .A1(n750), .A2(n735), .ZN(n105) );
endmodule


module FIR_Processor_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  CMPE32D1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  CMPE32D1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  CMPE32D1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  CMPE32D1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  CMPE32D1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  CMPE32D1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  CMPE32D1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  CMPE32D1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  CMPE32D1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  CMPE32D1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  CMPE32D1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  CMPE32D1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  CMPE32D1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  CMPE32D1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  CMPE32D1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  CMPE32D1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  CMPE32D1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  CMPE32D1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  CMPE32D1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  CMPE32D1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  CMPE32D1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  CMPE32D1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  CMPE32D1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  CMPE32D1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  CMPE32D1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  CMPE32D1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  CMPE32D1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  CMPE32D1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  CMPE32D1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  CMPE32D1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3D1 U1_31 ( .A1(A[31]), .A2(B[31]), .A3(carry[31]), .Z(SUM[31]) );
  AN2D0 U1 ( .A1(B[0]), .A2(A[0]), .Z(n1) );
  XOR2D1 U2 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module FIR_Processor ( rst_n, clk, sample_clk, sample_delay_in, coeficient, 
        coef_addr, dav, outp );
  input [15:0] sample_delay_in;
  input [15:0] coeficient;
  output [2:0] coef_addr;
  output [15:0] outp;
  input rst_n, clk, sample_clk;
  output dav;
  wire   CURRENT_STATE, NEXT_STATE, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45,
         N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59,
         N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N109,
         N110, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120,
         N121, N122, N123, N124, N125, N126, N127, N128, N129, N130, N131,
         N132, N133, N134, N135, N136, N137, N138, N139, N140, N176, N177,
         N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188,
         N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199,
         N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, n7,
         n8, n9, n10, n12, n13, n14, n15, n16, n18, n19, n20, n21, N99, N98,
         N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84,
         N83, N82, N81, N80, N79, N78, N77, N108, N107, N106, N105, N104, N103,
         N102, N101, N100, n1, n2, n3, n4, n5, n6, n11, n17, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31;
  wire   [31:0] counter;
  wire   [31:0] accumulator;

  IAO21D1 U39 ( .A1(n1), .A2(coef_addr[1]), .B(N208), .ZN(n9) );
  FIR_Processor_DW01_dec_0 sub_79 ( .A(counter), .SUM({N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, 
        N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9}) );
  FIR_Processor_DW_mult_uns_0 mult_115 ( .a(sample_delay_in), .b(coeficient), 
        .product({N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, 
        N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, 
        N84, N83, N82, N81, N80, N79, N78, N77}) );
  FIR_Processor_DW01_add_0 add_115 ( .A({N108, N107, N106, N105, N104, N103, 
        N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, 
        N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77}), .B(
        accumulator), .CI(1'b0), .SUM({N140, N139, N138, N137, N136, N135, 
        N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, 
        N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, 
        N110, N109}) );
  DFCNQD1 \accumulator_reg[31]  ( .D(N207), .CP(clk), .CDN(n24), .Q(
        accumulator[31]) );
  DFCNQD1 \accumulator_reg[30]  ( .D(N206), .CP(clk), .CDN(n24), .Q(
        accumulator[30]) );
  DFCNQD1 \accumulator_reg[29]  ( .D(N205), .CP(clk), .CDN(n25), .Q(
        accumulator[29]) );
  DFCNQD1 \accumulator_reg[28]  ( .D(N204), .CP(clk), .CDN(n25), .Q(
        accumulator[28]) );
  DFCNQD1 \accumulator_reg[27]  ( .D(N203), .CP(clk), .CDN(n25), .Q(
        accumulator[27]) );
  DFCNQD1 \accumulator_reg[26]  ( .D(N202), .CP(clk), .CDN(n25), .Q(
        accumulator[26]) );
  DFCNQD1 \accumulator_reg[25]  ( .D(N201), .CP(clk), .CDN(n25), .Q(
        accumulator[25]) );
  DFCNQD1 \accumulator_reg[24]  ( .D(N200), .CP(clk), .CDN(n25), .Q(
        accumulator[24]) );
  DFCNQD1 \accumulator_reg[23]  ( .D(N199), .CP(clk), .CDN(n25), .Q(
        accumulator[23]) );
  DFCNQD1 \accumulator_reg[22]  ( .D(N198), .CP(clk), .CDN(n25), .Q(
        accumulator[22]) );
  DFCNQD1 \accumulator_reg[21]  ( .D(N197), .CP(clk), .CDN(n25), .Q(
        accumulator[21]) );
  DFCNQD1 \accumulator_reg[20]  ( .D(N196), .CP(clk), .CDN(n25), .Q(
        accumulator[20]) );
  DFCNQD1 \counter_reg[31]  ( .D(N72), .CP(clk), .CDN(n24), .Q(counter[31]) );
  DFCNQD1 \counter_reg[27]  ( .D(N68), .CP(clk), .CDN(n24), .Q(counter[27]) );
  DFCNQD1 \counter_reg[29]  ( .D(N70), .CP(clk), .CDN(n24), .Q(counter[29]) );
  DFCNQD1 \counter_reg[25]  ( .D(N66), .CP(clk), .CDN(n23), .Q(counter[25]) );
  DFCNQD1 \counter_reg[26]  ( .D(N67), .CP(clk), .CDN(n24), .Q(counter[26]) );
  DFCNQD1 \counter_reg[28]  ( .D(N69), .CP(clk), .CDN(n24), .Q(counter[28]) );
  DFCNQD1 \counter_reg[30]  ( .D(N71), .CP(clk), .CDN(n24), .Q(counter[30]) );
  DFCNQD1 CURRENT_STATE_reg ( .D(NEXT_STATE), .CP(clk), .CDN(n24), .Q(
        CURRENT_STATE) );
  DFCNQD1 \accumulator_reg[19]  ( .D(N195), .CP(clk), .CDN(n25), .Q(
        accumulator[19]) );
  DFCNQD1 \accumulator_reg[18]  ( .D(N194), .CP(clk), .CDN(n26), .Q(
        accumulator[18]) );
  DFCNQD1 \accumulator_reg[17]  ( .D(N193), .CP(clk), .CDN(n26), .Q(
        accumulator[17]) );
  DFCNQD1 \accumulator_reg[16]  ( .D(N192), .CP(clk), .CDN(n26), .Q(
        accumulator[16]) );
  DFCNQD1 \accumulator_reg[15]  ( .D(N191), .CP(clk), .CDN(n26), .Q(
        accumulator[15]) );
  DFCNQD1 \accumulator_reg[14]  ( .D(N190), .CP(clk), .CDN(n26), .Q(
        accumulator[14]) );
  DFCNQD1 \accumulator_reg[13]  ( .D(N189), .CP(clk), .CDN(n26), .Q(
        accumulator[13]) );
  DFCNQD1 \accumulator_reg[12]  ( .D(N188), .CP(clk), .CDN(n26), .Q(
        accumulator[12]) );
  DFCNQD1 \accumulator_reg[11]  ( .D(N187), .CP(clk), .CDN(n26), .Q(
        accumulator[11]) );
  DFCNQD1 \accumulator_reg[10]  ( .D(N186), .CP(clk), .CDN(n26), .Q(
        accumulator[10]) );
  DFCNQD1 \accumulator_reg[9]  ( .D(N185), .CP(clk), .CDN(n26), .Q(
        accumulator[9]) );
  DFCNQD1 \accumulator_reg[8]  ( .D(N184), .CP(clk), .CDN(n25), .Q(
        accumulator[8]) );
  DFCNQD1 \accumulator_reg[7]  ( .D(N183), .CP(clk), .CDN(n26), .Q(
        accumulator[7]) );
  DFCNQD1 \accumulator_reg[6]  ( .D(N182), .CP(clk), .CDN(n26), .Q(
        accumulator[6]) );
  DFCNQD1 \accumulator_reg[5]  ( .D(N181), .CP(clk), .CDN(n27), .Q(
        accumulator[5]) );
  DFCNQD1 \accumulator_reg[4]  ( .D(N180), .CP(clk), .CDN(n27), .Q(
        accumulator[4]) );
  DFCNQD1 \counter_reg[16]  ( .D(N57), .CP(clk), .CDN(n23), .Q(counter[16]) );
  DFCNQD1 \counter_reg[23]  ( .D(N64), .CP(clk), .CDN(n23), .Q(counter[23]) );
  DFCNQD1 \counter_reg[15]  ( .D(N56), .CP(clk), .CDN(n23), .Q(counter[15]) );
  DFCNQD1 \counter_reg[19]  ( .D(N60), .CP(clk), .CDN(n23), .Q(counter[19]) );
  DFCNQD1 \counter_reg[22]  ( .D(N63), .CP(clk), .CDN(n23), .Q(counter[22]) );
  DFCNQD1 \counter_reg[14]  ( .D(N55), .CP(clk), .CDN(n23), .Q(counter[14]) );
  DFCNQD1 \counter_reg[18]  ( .D(N59), .CP(clk), .CDN(n23), .Q(counter[18]) );
  DFCNQD1 \counter_reg[21]  ( .D(N62), .CP(clk), .CDN(n23), .Q(counter[21]) );
  DFCNQD1 \counter_reg[17]  ( .D(N58), .CP(clk), .CDN(n23), .Q(counter[17]) );
  DFCNQD1 \counter_reg[20]  ( .D(N61), .CP(clk), .CDN(n23), .Q(counter[20]) );
  DFCNQD1 \counter_reg[24]  ( .D(N65), .CP(clk), .CDN(n23), .Q(counter[24]) );
  DFCNQD1 \accumulator_reg[3]  ( .D(N179), .CP(clk), .CDN(n27), .Q(
        accumulator[3]) );
  DFCNQD1 \accumulator_reg[2]  ( .D(N178), .CP(clk), .CDN(n27), .Q(
        accumulator[2]) );
  DFCNQD1 \accumulator_reg[1]  ( .D(N177), .CP(clk), .CDN(n27), .Q(
        accumulator[1]) );
  DFCNQD1 \counter_reg[12]  ( .D(N53), .CP(clk), .CDN(n22), .Q(counter[12]) );
  DFCNQD1 \counter_reg[8]  ( .D(N49), .CP(clk), .CDN(n22), .Q(counter[8]) );
  DFCNQD1 \counter_reg[6]  ( .D(N47), .CP(clk), .CDN(n22), .Q(counter[6]) );
  DFCNQD1 \counter_reg[13]  ( .D(N54), .CP(clk), .CDN(n22), .Q(counter[13]) );
  DFCNQD1 \counter_reg[9]  ( .D(N50), .CP(clk), .CDN(n22), .Q(counter[9]) );
  DFCNQD1 \counter_reg[7]  ( .D(N48), .CP(clk), .CDN(n22), .Q(counter[7]) );
  DFCNQD1 \accumulator_reg[0]  ( .D(N176), .CP(clk), .CDN(n27), .Q(
        accumulator[0]) );
  DFCNQD1 \counter_reg[10]  ( .D(N51), .CP(clk), .CDN(n22), .Q(counter[10]) );
  DFCNQD1 \counter_reg[11]  ( .D(N52), .CP(clk), .CDN(n22), .Q(counter[11]) );
  DFCNQD1 \coef_addr_wire_reg[2]  ( .D(N210), .CP(clk), .CDN(n24), .Q(
        coef_addr[2]) );
  DFCNQD1 \coef_addr_wire_reg[1]  ( .D(N209), .CP(clk), .CDN(n24), .Q(
        coef_addr[1]) );
  DFCNQD1 \counter_reg[1]  ( .D(N42), .CP(clk), .CDN(n22), .Q(counter[1]) );
  DFCNQD1 \counter_reg[5]  ( .D(N46), .CP(clk), .CDN(n22), .Q(counter[5]) );
  DFCNQD1 \counter_reg[4]  ( .D(N45), .CP(clk), .CDN(n22), .Q(counter[4]) );
  DFCNQD1 \counter_reg[3]  ( .D(N44), .CP(clk), .CDN(n22), .Q(counter[3]) );
  DFSND1 \counter_reg[0]  ( .D(N41), .CP(clk), .SDN(n27), .Q(counter[0]), .QN(
        n2) );
  DFSND1 \counter_reg[2]  ( .D(N43), .CP(clk), .SDN(n27), .Q(counter[2]) );
  DFCNQD1 \coef_addr_wire_reg[0]  ( .D(N208), .CP(clk), .CDN(n24), .Q(
        coef_addr[0]) );
  DFSND1 dav_wire_reg ( .D(n30), .CP(clk), .SDN(n27), .Q(dav) );
  EDFCNQD1 \outp_wire_reg[15]  ( .D(accumulator[15]), .E(n30), .CP(clk), .CDN(
        n27), .Q(outp[15]) );
  EDFCNQD1 \outp_wire_reg[14]  ( .D(accumulator[14]), .E(n30), .CP(clk), .CDN(
        n27), .Q(outp[14]) );
  EDFCNQD1 \outp_wire_reg[13]  ( .D(accumulator[13]), .E(n30), .CP(clk), .CDN(
        n28), .Q(outp[13]) );
  EDFCNQD1 \outp_wire_reg[12]  ( .D(accumulator[12]), .E(n30), .CP(clk), .CDN(
        n27), .Q(outp[12]) );
  EDFCNQD1 \outp_wire_reg[11]  ( .D(accumulator[11]), .E(n30), .CP(clk), .CDN(
        n27), .Q(outp[11]) );
  EDFCNQD1 \outp_wire_reg[10]  ( .D(accumulator[10]), .E(n30), .CP(clk), .CDN(
        n28), .Q(outp[10]) );
  EDFCNQD1 \outp_wire_reg[9]  ( .D(accumulator[9]), .E(n30), .CP(clk), .CDN(
        n28), .Q(outp[9]) );
  EDFCNQD1 \outp_wire_reg[8]  ( .D(accumulator[8]), .E(n30), .CP(clk), .CDN(
        n28), .Q(outp[8]) );
  EDFCNQD1 \outp_wire_reg[7]  ( .D(accumulator[7]), .E(n30), .CP(clk), .CDN(
        n28), .Q(outp[7]) );
  EDFCNQD1 \outp_wire_reg[6]  ( .D(accumulator[6]), .E(n30), .CP(clk), .CDN(
        n28), .Q(outp[6]) );
  EDFCNQD1 \outp_wire_reg[5]  ( .D(accumulator[5]), .E(n30), .CP(clk), .CDN(
        n28), .Q(outp[5]) );
  EDFCNQD1 \outp_wire_reg[4]  ( .D(accumulator[4]), .E(n30), .CP(clk), .CDN(
        n28), .Q(outp[4]) );
  EDFCNQD1 \outp_wire_reg[3]  ( .D(accumulator[3]), .E(n30), .CP(clk), .CDN(
        n28), .Q(outp[3]) );
  EDFCNQD1 \outp_wire_reg[2]  ( .D(accumulator[2]), .E(n30), .CP(clk), .CDN(
        n28), .Q(outp[2]) );
  EDFCNQD1 \outp_wire_reg[1]  ( .D(accumulator[1]), .E(n30), .CP(clk), .CDN(
        n28), .Q(outp[1]) );
  EDFCNQD1 \outp_wire_reg[0]  ( .D(accumulator[0]), .E(n30), .CP(clk), .CDN(
        n28), .Q(outp[0]) );
  AO21D1 U3 ( .A1(n29), .A2(counter[2]), .B(n30), .Z(n1) );
  BUFFD0 U4 ( .I(n17), .Z(n28) );
  INVD1 U5 ( .I(sample_clk), .ZN(n5) );
  AN2D0 U6 ( .A1(N38), .A2(n5), .Z(N70) );
  AN2D0 U7 ( .A1(N36), .A2(n5), .Z(N68) );
  AN2D0 U8 ( .A1(N128), .A2(n4), .Z(N195) );
  AN2D0 U9 ( .A1(N129), .A2(n4), .Z(N196) );
  AN2D0 U10 ( .A1(N130), .A2(n4), .Z(N197) );
  AN2D0 U11 ( .A1(N131), .A2(n4), .Z(N198) );
  AN2D0 U12 ( .A1(N132), .A2(n4), .Z(N199) );
  AN2D0 U13 ( .A1(N133), .A2(n4), .Z(N200) );
  AN2D0 U14 ( .A1(N134), .A2(n4), .Z(N201) );
  AN2D0 U15 ( .A1(N135), .A2(n4), .Z(N202) );
  AN2D0 U16 ( .A1(N136), .A2(n4), .Z(N203) );
  AN2D0 U17 ( .A1(N137), .A2(n4), .Z(N204) );
  AN2D0 U18 ( .A1(N138), .A2(n4), .Z(N205) );
  AN2D0 U19 ( .A1(N139), .A2(n4), .Z(N206) );
  AN2D0 U20 ( .A1(N17), .A2(n5), .Z(N49) );
  AN2D0 U21 ( .A1(N21), .A2(n5), .Z(N53) );
  AN2D0 U22 ( .A1(N19), .A2(n5), .Z(N51) );
  AN2D0 U23 ( .A1(N112), .A2(n4), .Z(N179) );
  AN2D0 U24 ( .A1(N113), .A2(n4), .Z(N180) );
  AN2D0 U25 ( .A1(N114), .A2(n4), .Z(N181) );
  AN2D0 U26 ( .A1(N115), .A2(n4), .Z(N182) );
  AN2D0 U27 ( .A1(N116), .A2(n4), .Z(N183) );
  AN2D0 U28 ( .A1(N117), .A2(n4), .Z(N184) );
  AN2D0 U29 ( .A1(N118), .A2(n4), .Z(N185) );
  AN2D0 U30 ( .A1(N119), .A2(n4), .Z(N186) );
  AN2D0 U31 ( .A1(N120), .A2(n4), .Z(N187) );
  AN2D0 U32 ( .A1(N121), .A2(n4), .Z(N188) );
  AN2D0 U33 ( .A1(N122), .A2(n4), .Z(N189) );
  AN2D0 U34 ( .A1(N123), .A2(n4), .Z(N190) );
  AN2D0 U35 ( .A1(N124), .A2(n4), .Z(N191) );
  AN2D0 U36 ( .A1(N125), .A2(n4), .Z(N192) );
  AN2D0 U37 ( .A1(N126), .A2(n4), .Z(N193) );
  AN2D0 U38 ( .A1(N127), .A2(n4), .Z(N194) );
  INVD1 U40 ( .I(n1), .ZN(n4) );
  AN2D0 U41 ( .A1(N111), .A2(n4), .Z(N178) );
  AN2D0 U42 ( .A1(N110), .A2(n4), .Z(N177) );
  BUFFD0 U43 ( .I(n11), .Z(n27) );
  BUFFD0 U44 ( .I(n11), .Z(n26) );
  BUFFD0 U45 ( .I(n11), .Z(n25) );
  BUFFD0 U46 ( .I(n6), .Z(n24) );
  BUFFD0 U47 ( .I(n6), .Z(n23) );
  BUFFD0 U48 ( .I(n6), .Z(n22) );
  AN2D0 U49 ( .A1(N140), .A2(n4), .Z(N207) );
  AN2D0 U50 ( .A1(N40), .A2(n5), .Z(N72) );
  AN2D0 U51 ( .A1(N39), .A2(n5), .Z(N71) );
  AN2D0 U52 ( .A1(N37), .A2(n5), .Z(N69) );
  AN2D0 U53 ( .A1(N35), .A2(n5), .Z(N67) );
  AN2D0 U54 ( .A1(N34), .A2(n5), .Z(N66) );
  AN2D0 U55 ( .A1(N33), .A2(n5), .Z(N65) );
  AN2D0 U56 ( .A1(N32), .A2(n5), .Z(N64) );
  AN2D0 U57 ( .A1(N31), .A2(n5), .Z(N63) );
  AN2D0 U58 ( .A1(N30), .A2(n5), .Z(N62) );
  AN2D0 U59 ( .A1(N29), .A2(n5), .Z(N61) );
  AN2D0 U60 ( .A1(N28), .A2(n5), .Z(N60) );
  AN2D0 U61 ( .A1(N27), .A2(n5), .Z(N59) );
  AN2D0 U62 ( .A1(N26), .A2(n5), .Z(N58) );
  AN2D0 U63 ( .A1(N20), .A2(n5), .Z(N52) );
  AN2D0 U64 ( .A1(N25), .A2(n5), .Z(N57) );
  AN2D0 U65 ( .A1(N24), .A2(n5), .Z(N56) );
  AN2D0 U66 ( .A1(N23), .A2(n5), .Z(N55) );
  AN2D0 U67 ( .A1(N22), .A2(n5), .Z(N54) );
  AN2D0 U68 ( .A1(N18), .A2(n5), .Z(N50) );
  NR4D0 U69 ( .A1(counter[26]), .A2(counter[25]), .A3(counter[24]), .A4(
        counter[23]), .ZN(n18) );
  NR4D0 U70 ( .A1(counter[9]), .A2(counter[8]), .A3(counter[7]), .A4(
        counter[6]), .ZN(n21) );
  NR4D0 U71 ( .A1(counter[5]), .A2(counter[4]), .A3(counter[3]), .A4(
        counter[31]), .ZN(n20) );
  NR4D0 U72 ( .A1(counter[30]), .A2(counter[29]), .A3(counter[28]), .A4(
        counter[27]), .ZN(n19) );
  IND2D1 U73 ( .A1(N11), .B1(n5), .ZN(N43) );
  OAI22D0 U74 ( .A1(CURRENT_STATE), .A2(n5), .B1(n30), .B2(n7), .ZN(NEXT_STATE) );
  NR2D1 U75 ( .A1(counter[2]), .A2(n8), .ZN(n7) );
  OAI21D0 U76 ( .A1(n9), .A2(n31), .B(n10), .ZN(N210) );
  ND4D1 U77 ( .A1(coef_addr[1]), .A2(coef_addr[0]), .A3(n4), .A4(n31), .ZN(n10) );
  INVD1 U78 ( .I(coef_addr[2]), .ZN(n31) );
  INVD1 U79 ( .I(n8), .ZN(n29) );
  INVD1 U80 ( .I(CURRENT_STATE), .ZN(n30) );
  NR4D0 U81 ( .A1(n2), .A2(n3), .A3(counter[11]), .A4(counter[10]), .ZN(n15)
         );
  OR4D1 U82 ( .A1(counter[15]), .A2(counter[14]), .A3(counter[13]), .A4(
        counter[12]), .Z(n3) );
  IND4D1 U83 ( .A1(n13), .B1(n14), .B2(n15), .B3(n16), .ZN(n8) );
  NR4D0 U84 ( .A1(counter[19]), .A2(counter[18]), .A3(counter[17]), .A4(
        counter[16]), .ZN(n16) );
  NR4D0 U85 ( .A1(counter[22]), .A2(counter[21]), .A3(counter[20]), .A4(
        counter[1]), .ZN(n14) );
  ND4D1 U86 ( .A1(n18), .A2(n19), .A3(n20), .A4(n21), .ZN(n13) );
  NR2D1 U87 ( .A1(n1), .A2(coef_addr[0]), .ZN(N208) );
  AN2D0 U88 ( .A1(N14), .A2(n5), .Z(N46) );
  AN2D0 U89 ( .A1(N12), .A2(n5), .Z(N44) );
  AN2D0 U90 ( .A1(N16), .A2(n5), .Z(N48) );
  NR2D1 U91 ( .A1(n12), .A2(n1), .ZN(N209) );
  XNR2D1 U92 ( .A1(coef_addr[1]), .A2(coef_addr[0]), .ZN(n12) );
  AN2D0 U93 ( .A1(N109), .A2(n4), .Z(N176) );
  AN2D0 U94 ( .A1(N15), .A2(n5), .Z(N47) );
  AN2D0 U95 ( .A1(N13), .A2(n5), .Z(N45) );
  AN2D0 U96 ( .A1(N10), .A2(n5), .Z(N42) );
  IND2D1 U97 ( .A1(N9), .B1(n5), .ZN(N41) );
  BUFFD0 U98 ( .I(rst_n), .Z(n17) );
  BUFFD0 U99 ( .I(rst_n), .Z(n6) );
  BUFFD0 U100 ( .I(rst_n), .Z(n11) );
endmodule


module ROM_Process ( address, coeficient_out );
  input [2:0] address;
  output [15:0] coeficient_out;
  wire   \address[2] , n1, n2;
  assign coeficient_out[4] = 1'b0;
  assign coeficient_out[5] = 1'b0;
  assign coeficient_out[6] = 1'b0;
  assign coeficient_out[7] = 1'b0;
  assign coeficient_out[8] = 1'b0;
  assign coeficient_out[9] = 1'b0;
  assign coeficient_out[10] = 1'b0;
  assign coeficient_out[11] = 1'b0;
  assign coeficient_out[12] = 1'b0;
  assign coeficient_out[13] = 1'b0;
  assign coeficient_out[14] = 1'b0;
  assign coeficient_out[15] = 1'b0;
  assign coeficient_out[3] = \address[2] ;
  assign \address[2]  = address[2];

  NR2D1 U3 ( .A1(coeficient_out[1]), .A2(n1), .ZN(coeficient_out[2]) );
  XNR2D1 U4 ( .A1(address[1]), .A2(n1), .ZN(coeficient_out[1]) );
  INVD1 U5 ( .I(address[0]), .ZN(n1) );
  AOI21D0 U6 ( .A1(\address[2] ), .A2(n2), .B(address[0]), .ZN(
        coeficient_out[0]) );
  INVD1 U7 ( .I(address[1]), .ZN(n2) );
endmodule


module FIR_Toplevel ( rst_n, clk, sample_clk, sample, dav, outp );
  input [15:0] sample;
  output [15:0] outp;
  input rst_n, clk, sample_clk;
  output dav;

  wire   [15:0] sample_out_wire;
  wire   [15:0] coeficient_out_wire;
  wire   [2:0] coef_addr_wire;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11;

  Delayline_CB U_delayline ( .rst_n(rst_n), .clk(clk), .sample_clk(sample_clk), 
        .sample(sample), .sample_out(sample_out_wire) );
  FIR_Processor u_FIRP ( .rst_n(rst_n), .clk(clk), .sample_clk(sample_clk), 
        .sample_delay_in(sample_out_wire), .coeficient({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        coeficient_out_wire[3:0]}), .coef_addr(coef_addr_wire), .dav(dav), 
        .outp(outp) );
  ROM_Process u_ROM ( .address(coef_addr_wire), .coeficient_out({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        coeficient_out_wire[3:0]}) );
endmodule

