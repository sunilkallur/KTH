module add_6_100(A, B, Z);
    input [5 : 0] A;
    input [5 : 0] B;
    output [5 : 0] Z;

    assign Z = A + B;
endmodule
